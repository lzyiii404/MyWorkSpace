//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_194_assert(
  input  [3:0]  _EVAL_1,
  input         _EVAL_4,
  input  [6:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_71,
  input         _EVAL_114,
  input         _EVAL_59,
  input  [31:0] _EVAL_81,
  input         _EVAL_98,
  input         _EVAL_56,
  input         _EVAL_139,
  input         _EVAL_25,
  input         _EVAL_122,
  input         _EVAL_117,
  input         _EVAL_49,
  input         _EVAL_66,
  input         _EVAL_129,
  input         _EVAL_74,
  input         _EVAL_130,
  input         _EVAL_133,
  input         _EVAL_107,
  input         _EVAL_50,
  input         _EVAL_27
);
  wire  TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire [2:0] TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire [3:0] TLMonitor__EVAL_4;
  wire [6:0] TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  _EVAL_61;
  wire  _EVAL_83;
  wire  _EVAL_106;
  wire  _EVAL_54;
  wire  _EVAL_20;
  wire  _EVAL_51;
  wire  _EVAL_44;
  wire [11:0] _EVAL_72;
  wire  _EVAL_46;
  wire  _EVAL_108;
  wire  _EVAL_100;
  wire  _EVAL_132;
  wire  _EVAL_95;
  wire  _EVAL_70;
  wire  _EVAL_101;
  wire  _EVAL_140;
  wire  _EVAL_42;
  wire  _EVAL_69;
  wire [8:0] _EVAL_92;
  wire  _EVAL_24;
  wire  _EVAL_93;
  wire  _EVAL_89;
  wire  _EVAL_105;
  wire  _EVAL_136;
  wire  _EVAL_39;
  wire  _EVAL_79;
  wire  _EVAL_115;
  wire  _EVAL_48;
  wire  _EVAL_128;
  wire  _EVAL_116;
  wire  _EVAL_23;
  wire  _EVAL_103;
  SiFive__EVAL_191_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8)
  );
  assign _EVAL_61 = _EVAL_71 & _EVAL_114;
  assign _EVAL_83 = _EVAL_61 & _EVAL_59;
  assign _EVAL_106 = _EVAL_83 & _EVAL_98;
  assign _EVAL_54 = _EVAL_83 & _EVAL_25;
  assign _EVAL_20 = _EVAL_83 & _EVAL_122;
  assign _EVAL_51 = _EVAL_81[29];
  assign _EVAL_44 = _EVAL_56 & _EVAL_51;
  assign _EVAL_72 = _EVAL_81[15:4];
  assign _EVAL_46 = _EVAL_72 == 12'hfff;
  assign _EVAL_108 = _EVAL_56 & _EVAL_46;
  assign _EVAL_100 = _EVAL_81[26];
  assign _EVAL_132 = _EVAL_83 & _EVAL_100;
  assign _EVAL_95 = _EVAL_81[16];
  assign _EVAL_70 = _EVAL_83 & _EVAL_95;
  assign _EVAL_101 = _EVAL_72 != 12'h0;
  assign _EVAL_140 = _EVAL_83 & _EVAL_101;
  assign _EVAL_42 = _EVAL_81[27];
  assign _EVAL_69 = _EVAL_83 & _EVAL_42;
  assign _EVAL_92 = _EVAL_81[25:17];
  assign _EVAL_24 = _EVAL_92 == 9'h1ff;
  assign _EVAL_93 = _EVAL_56 & _EVAL_100;
  assign _EVAL_89 = _EVAL_83 & _EVAL_130;
  assign _EVAL_105 = _EVAL_83 & _EVAL_51;
  assign _EVAL_136 = _EVAL_83 & _EVAL_74;
  assign _EVAL_39 = _EVAL_83 & _EVAL_66;
  assign _EVAL_79 = _EVAL_92 != 9'h0;
  assign _EVAL_115 = _EVAL_56 & _EVAL_95;
  assign _EVAL_48 = _EVAL_83 & _EVAL_49;
  assign _EVAL_128 = _EVAL_83 & _EVAL_79;
  assign _EVAL_116 = _EVAL_4 == 1'h0;
  assign _EVAL_23 = _EVAL_56 & _EVAL_42;
  assign _EVAL_103 = _EVAL_56 & _EVAL_24;
  assign TLMonitor__EVAL_4 = _EVAL_1;
  assign TLMonitor__EVAL_6 = _EVAL_13;
  assign TLMonitor__EVAL_3 = _EVAL_9;
  assign TLMonitor__EVAL_0 = _EVAL_14;
  assign TLMonitor__EVAL_8 = _EVAL_13;
  assign TLMonitor__EVAL_7 = _EVAL_9;
  assign TLMonitor__EVAL_5 = _EVAL_8;
  assign TLMonitor__EVAL = _EVAL_4;
  assign TLMonitor__EVAL_2 = {{2'd0}, _EVAL_114};
  assign TLMonitor__EVAL_1 = _EVAL_15;
  always @(posedge _EVAL_14) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f62378dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b7373ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e585bfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15caf87e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bfc75b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd8f979e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53661116)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(139303cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbaf213a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f291f85a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6918a3ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c4bac4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(210fe89e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5d69497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaf5be21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a84dc116)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ecd8080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99f7ad2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(368a3af5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48c4c0ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c2be1c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad56e30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98d393d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e512a2e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d839b96e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f1aec64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(468ebe99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b24dc15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(399a8720)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3482d9eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e739463d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e7e400e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
