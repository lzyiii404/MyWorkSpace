//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_225_assert(
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_9,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [31:0] _EVAL_17,
  input         _EVAL_19,
  input  [3:0]  _EVAL_20,
  input  [31:0] _EVAL_22,
  input         _EVAL_23,
  input  [3:0]  _EVAL_26,
  input         _EVAL_28,
  input  [2:0]  _EVAL_29,
  input         _EVAL_44,
  input  [3:0]  _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_50,
  input         _EVAL_51,
  input  [2:0]  _EVAL_52,
  input         _EVAL_53,
  input  [2:0]  _EVAL_56,
  input         _EVAL_59,
  input         _EVAL_60,
  input  [2:0]  _EVAL_61,
  input         _EVAL_67,
  input  [1:0]  _EVAL_68,
  input  [31:0] _EVAL_70,
  input         _EVAL_71,
  input  [2:0]  _EVAL_74,
  input         _EVAL_75,
  input  [1:0]  _EVAL_76,
  input  [7:0]  _EVAL_77,
  input  [2:0]  _EVAL_79,
  input         _EVAL_80,
  input         _EVAL_81,
  input  [31:0] _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  input  [1:0]  _EVAL_98,
  input         _EVAL_133,
  input         _EVAL_146,
  input         _EVAL_121,
  input         _EVAL_94,
  input         _EVAL_87,
  input         _EVAL_118
);
  wire  TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [1:0] TLMonitor__EVAL_7;
  wire [31:0] TLMonitor__EVAL_8;
  wire [3:0] TLMonitor__EVAL_9;
  wire [2:0] TLMonitor__EVAL_10;
  wire  TLMonitor_1__EVAL;
  wire [2:0] TLMonitor_1__EVAL_0;
  wire  TLMonitor_1__EVAL_1;
  wire [1:0] TLMonitor_1__EVAL_2;
  wire [7:0] TLMonitor_1__EVAL_3;
  wire [3:0] TLMonitor_1__EVAL_4;
  wire  TLMonitor_1__EVAL_5;
  wire [2:0] TLMonitor_1__EVAL_6;
  wire [2:0] TLMonitor_1__EVAL_7;
  wire [2:0] TLMonitor_1__EVAL_8;
  wire  TLMonitor_1__EVAL_9;
  wire  TLMonitor_1__EVAL_10;
  wire  TLMonitor_1__EVAL_11;
  wire [2:0] TLMonitor_1__EVAL_12;
  wire  TLMonitor_1__EVAL_13;
  wire [1:0] TLMonitor_1__EVAL_14;
  wire [2:0] TLMonitor_1__EVAL_15;
  wire  TLMonitor_1__EVAL_16;
  wire  TLMonitor_1__EVAL_17;
  wire  TLMonitor_1__EVAL_18;
  wire  TLMonitor_1__EVAL_19;
  wire [3:0] TLMonitor_1__EVAL_20;
  wire [31:0] TLMonitor_1__EVAL_21;
  wire  TLMonitor_1__EVAL_22;
  wire  TLMonitor_1__EVAL_23;
  wire [31:0] TLMonitor_1__EVAL_24;
  wire [31:0] TLMonitor_1__EVAL_25;
  wire  TLMonitor_1__EVAL_26;
  wire  TLMonitor_1__EVAL_27;
  wire [3:0] TLMonitor_1__EVAL_28;
  wire [2:0] TLMonitor_1__EVAL_29;
  wire  TLMonitor_1__EVAL_30;
  wire  TLMonitor_1__EVAL_31;
  wire  TLMonitor_1__EVAL_32;
  wire [2:0] TLMonitor_1__EVAL_33;
  wire  _EVAL_114;
  wire  _EVAL_141;
  wire  _EVAL_95;
  wire  _EVAL_122;
  wire  _EVAL_111;
  wire  _EVAL_130;
  wire  _EVAL_109;
  wire  _EVAL_147;
  wire  _EVAL_138;
  wire  _EVAL_101;
  wire  _EVAL_124;
  wire  _EVAL_145;
  wire  _EVAL_120;
  SiFive__EVAL_223_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10)
  );
  SiFive__EVAL_224_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14),
    ._EVAL_15(TLMonitor_1__EVAL_15),
    ._EVAL_16(TLMonitor_1__EVAL_16),
    ._EVAL_17(TLMonitor_1__EVAL_17),
    ._EVAL_18(TLMonitor_1__EVAL_18),
    ._EVAL_19(TLMonitor_1__EVAL_19),
    ._EVAL_20(TLMonitor_1__EVAL_20),
    ._EVAL_21(TLMonitor_1__EVAL_21),
    ._EVAL_22(TLMonitor_1__EVAL_22),
    ._EVAL_23(TLMonitor_1__EVAL_23),
    ._EVAL_24(TLMonitor_1__EVAL_24),
    ._EVAL_25(TLMonitor_1__EVAL_25),
    ._EVAL_26(TLMonitor_1__EVAL_26),
    ._EVAL_27(TLMonitor_1__EVAL_27),
    ._EVAL_28(TLMonitor_1__EVAL_28),
    ._EVAL_29(TLMonitor_1__EVAL_29),
    ._EVAL_30(TLMonitor_1__EVAL_30),
    ._EVAL_31(TLMonitor_1__EVAL_31),
    ._EVAL_32(TLMonitor_1__EVAL_32),
    ._EVAL_33(TLMonitor_1__EVAL_33)
  );
  assign _EVAL_114 = _EVAL_121 == 1'h0;
  assign _EVAL_141 = _EVAL_133 == 1'h0;
  assign _EVAL_95 = _EVAL_114 | _EVAL_141;
  assign _EVAL_122 = _EVAL_95 | _EVAL_83;
  assign _EVAL_111 = _EVAL_122 == 1'h0;
  assign _EVAL_130 = _EVAL_121 | _EVAL_133;
  assign _EVAL_109 = _EVAL_98 == _EVAL_98;
  assign _EVAL_147 = _EVAL_84 == 1'h0;
  assign _EVAL_138 = _EVAL_147 | _EVAL_130;
  assign _EVAL_101 = _EVAL_138 | _EVAL_83;
  assign _EVAL_124 = _EVAL_101 == 1'h0;
  assign _EVAL_145 = _EVAL_109 | _EVAL_83;
  assign _EVAL_120 = _EVAL_145 == 1'h0;
  assign TLMonitor__EVAL_4 = _EVAL_60;
  assign TLMonitor_1__EVAL_23 = _EVAL_47;
  assign TLMonitor__EVAL_6 = _EVAL_51 & _EVAL_146;
  assign TLMonitor_1__EVAL_1 = _EVAL_59;
  assign TLMonitor_1__EVAL_21 = _EVAL_22;
  assign TLMonitor_1__EVAL_33 = _EVAL_79;
  assign TLMonitor_1__EVAL_6 = _EVAL_56;
  assign TLMonitor__EVAL_0 = _EVAL_75;
  assign TLMonitor__EVAL_9 = _EVAL_26;
  assign TLMonitor_1__EVAL_16 = _EVAL_13;
  assign TLMonitor_1__EVAL_3 = _EVAL_77;
  assign TLMonitor_1__EVAL_10 = _EVAL_4;
  assign TLMonitor_1__EVAL_26 = _EVAL_51 & _EVAL_87;
  assign TLMonitor_1__EVAL_29 = _EVAL_74;
  assign TLMonitor_1__EVAL_13 = _EVAL_19;
  assign TLMonitor__EVAL = _EVAL_47;
  assign TLMonitor_1__EVAL_15 = _EVAL_61;
  assign TLMonitor_1__EVAL_9 = _EVAL_44;
  assign TLMonitor_1__EVAL_30 = _EVAL_23;
  assign TLMonitor_1__EVAL_19 = _EVAL_75;
  assign TLMonitor_1__EVAL_4 = _EVAL_20;
  assign TLMonitor_1__EVAL_22 = _EVAL_71 & _EVAL_94;
  assign TLMonitor_1__EVAL_20 = _EVAL_26;
  assign TLMonitor_1__EVAL_25 = _EVAL_70;
  assign TLMonitor_1__EVAL_7 = _EVAL_29;
  assign TLMonitor_1__EVAL_11 = _EVAL_28;
  assign TLMonitor_1__EVAL_14 = _EVAL_76;
  assign TLMonitor__EVAL_3 = _EVAL_80;
  assign TLMonitor_1__EVAL_31 = _EVAL_81;
  assign TLMonitor__EVAL_2 = _EVAL_83;
  assign TLMonitor_1__EVAL_5 = _EVAL_83;
  assign TLMonitor__EVAL_1 = _EVAL_13;
  assign TLMonitor__EVAL_5 = _EVAL_71 & _EVAL_118;
  assign TLMonitor__EVAL_10 = _EVAL_29;
  assign TLMonitor__EVAL_8 = _EVAL_82;
  assign TLMonitor_1__EVAL_17 = _EVAL_53;
  assign TLMonitor_1__EVAL_2 = _EVAL_68;
  assign TLMonitor_1__EVAL_12 = _EVAL_3;
  assign TLMonitor_1__EVAL_24 = _EVAL_17;
  assign TLMonitor_1__EVAL_32 = _EVAL_50;
  assign TLMonitor_1__EVAL_18 = _EVAL_67;
  assign TLMonitor_1__EVAL_0 = _EVAL_46[2:0];
  assign TLMonitor__EVAL_7 = _EVAL_76;
  assign TLMonitor_1__EVAL = _EVAL_80;
  assign TLMonitor_1__EVAL_28 = _EVAL_14;
  assign TLMonitor_1__EVAL_27 = _EVAL_9;
  assign TLMonitor_1__EVAL_8 = _EVAL_52;
  always @(posedge _EVAL_80) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a924c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883ce8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0bb131)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
