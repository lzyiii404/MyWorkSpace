//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_310(
  output [31:0] _EVAL,
  input         _EVAL_0,
  output [31:0] _EVAL_1,
  input         _EVAL_2,
  output [63:0] _EVAL_3,
  output [2:0]  _EVAL_4,
  output [6:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  output [1:0]  _EVAL_10,
  output [3:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  output        _EVAL_13,
  input  [1:0]  _EVAL_14,
  output        _EVAL_15,
  output [7:0]  _EVAL_16,
  output        _EVAL_17,
  output [3:0]  _EVAL_18,
  input  [1:0]  _EVAL_19,
  output        _EVAL_20,
  input  [1:0]  _EVAL_21,
  input  [31:0] _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  output [7:0]  _EVAL_25,
  input  [31:0] _EVAL_26,
  output [31:0] _EVAL_27,
  input  [2:0]  _EVAL_28,
  output [3:0]  _EVAL_29,
  input  [1:0]  _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [2:0]  _EVAL_33,
  output [2:0]  _EVAL_34,
  output        _EVAL_35,
  input  [2:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  input  [31:0] _EVAL_38,
  input  [31:0] _EVAL_39,
  output [2:0]  _EVAL_40,
  input  [3:0]  _EVAL_41,
  input         _EVAL_42,
  output [1:0]  _EVAL_43,
  output        _EVAL_44,
  input  [63:0] _EVAL_45,
  output [3:0]  _EVAL_46,
  input         _EVAL_47,
  input  [6:0]  _EVAL_48,
  output [31:0] _EVAL_49,
  input  [31:0] _EVAL_50,
  input  [1:0]  _EVAL_51,
  output [1:0]  _EVAL_52,
  input         _EVAL_53,
  input  [1:0]  _EVAL_54,
  input  [2:0]  _EVAL_55,
  output [1:0]  _EVAL_56,
  output [3:0]  _EVAL_57,
  output [2:0]  _EVAL_58,
  input  [6:0]  _EVAL_59,
  output [1:0]  _EVAL_60,
  input  [1:0]  _EVAL_61,
  output [3:0]  _EVAL_62,
  input  [3:0]  _EVAL_63,
  input         _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_68,
  output        _EVAL_69,
  input  [1:0]  _EVAL_70,
  output [1:0]  _EVAL_71,
  input         _EVAL_72,
  output [2:0]  _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  output        _EVAL_76,
  output [2:0]  _EVAL_77,
  input  [63:0] _EVAL_78,
  output [2:0]  _EVAL_79,
  input         _EVAL_80,
  output [1:0]  _EVAL_81,
  output [31:0] _EVAL_82,
  input         _EVAL_83,
  input  [2:0]  _EVAL_84,
  output [6:0]  _EVAL_85,
  input  [1:0]  _EVAL_86,
  output        _EVAL_87,
  output [31:0] _EVAL_88,
  input         _EVAL_89,
  input  [24:0] _EVAL_90,
  input  [3:0]  _EVAL_91,
  output        _EVAL_92,
  output [3:0]  _EVAL_93,
  input  [2:0]  _EVAL_94,
  output        _EVAL_95,
  output [2:0]  _EVAL_96,
  output [2:0]  _EVAL_97,
  input  [24:0] _EVAL_98,
  output [3:0]  _EVAL_99,
  input         _EVAL_100,
  input         _EVAL_101,
  input         _EVAL_102,
  output [63:0] _EVAL_103,
  input  [3:0]  _EVAL_104,
  output        _EVAL_105,
  output [63:0] _EVAL_106,
  input  [3:0]  _EVAL_107,
  output [1:0]  _EVAL_108,
  output        _EVAL_109,
  output [1:0]  _EVAL_110,
  input  [1:0]  _EVAL_111,
  input         _EVAL_112,
  output        _EVAL_113,
  output [2:0]  _EVAL_114,
  input  [2:0]  _EVAL_115,
  output [63:0] _EVAL_116,
  output        _EVAL_117,
  output        _EVAL_118
);
  wire  fragmenter_1__EVAL;
  wire  fragmenter_1__EVAL_0;
  wire [1:0] fragmenter_1__EVAL_1;
  wire  fragmenter_1__EVAL_2;
  wire  fragmenter_1__EVAL_3;
  wire [7:0] fragmenter_1__EVAL_4;
  wire [2:0] fragmenter_1__EVAL_5;
  wire [2:0] fragmenter_1__EVAL_6;
  wire  fragmenter_1__EVAL_7;
  wire  fragmenter_1__EVAL_8;
  wire [3:0] fragmenter_1__EVAL_9;
  wire [31:0] fragmenter_1__EVAL_10;
  wire [24:0] fragmenter_1__EVAL_11;
  wire [2:0] fragmenter_1__EVAL_12;
  wire [2:0] fragmenter_1__EVAL_13;
  wire [31:0] fragmenter_1__EVAL_14;
  wire  fragmenter_1__EVAL_15;
  wire  fragmenter_1__EVAL_16;
  wire [3:0] fragmenter_1__EVAL_17;
  wire [7:0] fragmenter_1__EVAL_18;
  wire [31:0] fragmenter_1__EVAL_19;
  wire  fragmenter_1__EVAL_20;
  wire [2:0] fragmenter_1__EVAL_21;
  wire [1:0] fragmenter_1__EVAL_22;
  wire [31:0] fragmenter_1__EVAL_23;
  wire  fragmenter_1__EVAL_24;
  wire [24:0] fragmenter_1__EVAL_25;
  wire [2:0] fragmenter_1__EVAL_26;
  wire  fragmenter_1__EVAL_27;
  wire [12:0] fragmenter_1__EVAL_28;
  wire [2:0] fragmenter_1__EVAL_29;
  wire [12:0] fragmenter_1__EVAL_30;
  wire [2:0] fragmenter_1__EVAL_31;
  wire  fragmenter_1__EVAL_32;
  wire  dls__EVAL;
  wire [1:0] dls__EVAL_0;
  wire  dls__EVAL_1;
  wire [1:0] dls__EVAL_2;
  wire  dls__EVAL_3;
  wire [2:0] dls__EVAL_4;
  wire [3:0] dls__EVAL_5;
  wire  dls__EVAL_6;
  wire [12:0] dls__EVAL_7;
  wire  dls__EVAL_8;
  wire [2:0] dls__EVAL_9;
  wire [31:0] dls__EVAL_10;
  wire [24:0] dls__EVAL_11;
  wire [12:0] dls__EVAL_12;
  wire  dls__EVAL_13;
  wire [31:0] dls__EVAL_14;
  wire  dls__EVAL_15;
  wire [2:0] dls__EVAL_16;
  wire [2:0] widget__EVAL;
  wire [63:0] widget__EVAL_0;
  wire  widget__EVAL_1;
  wire [2:0] widget__EVAL_2;
  wire [6:0] widget__EVAL_3;
  wire [24:0] widget__EVAL_4;
  wire [2:0] widget__EVAL_5;
  wire [7:0] widget__EVAL_6;
  wire [2:0] widget__EVAL_7;
  wire  widget__EVAL_8;
  wire  widget__EVAL_9;
  wire  widget__EVAL_10;
  wire  widget__EVAL_11;
  wire  widget__EVAL_12;
  wire [2:0] widget__EVAL_13;
  wire [24:0] widget__EVAL_14;
  wire [6:0] widget__EVAL_15;
  wire [2:0] widget__EVAL_16;
  wire [3:0] widget__EVAL_17;
  wire [6:0] widget__EVAL_18;
  wire  widget__EVAL_19;
  wire  widget__EVAL_20;
  wire [6:0] widget__EVAL_21;
  wire [2:0] widget__EVAL_22;
  wire [63:0] widget__EVAL_23;
  wire [31:0] widget__EVAL_24;
  wire [2:0] widget__EVAL_25;
  wire  widget__EVAL_26;
  wire  widget__EVAL_27;
  wire [31:0] widget__EVAL_28;
  wire  dcache__EVAL;
  wire  dcache__EVAL_0;
  wire  dcache__EVAL_1;
  wire [29:0] dcache__EVAL_2;
  wire  dcache__EVAL_3;
  wire  dcache__EVAL_4;
  wire [2:0] dcache__EVAL_5;
  wire  dcache__EVAL_6;
  wire  dcache__EVAL_7;
  wire [31:0] dcache__EVAL_8;
  wire  dcache__EVAL_9;
  wire  dcache__EVAL_10;
  wire  dcache__EVAL_11;
  wire  dcache__EVAL_12;
  wire  dcache__EVAL_13;
  wire  dcache__EVAL_14;
  wire  dcache__EVAL_15;
  wire  dcache__EVAL_16;
  wire [5:0] dcache__EVAL_17;
  wire  dcache__EVAL_18;
  wire [29:0] dcache__EVAL_19;
  wire [31:0] dcache__EVAL_20;
  wire  dcache__EVAL_21;
  wire [31:0] dcache__EVAL_22;
  wire  dcache__EVAL_23;
  wire  dcache__EVAL_24;
  wire  dcache__EVAL_25;
  wire [29:0] dcache__EVAL_26;
  wire  dcache__EVAL_27;
  wire [29:0] dcache__EVAL_28;
  wire  dcache__EVAL_29;
  wire [2:0] dcache__EVAL_30;
  wire  dcache__EVAL_31;
  wire  dcache__EVAL_32;
  wire  dcache__EVAL_33;
  wire [1:0] dcache__EVAL_34;
  wire  dcache__EVAL_35;
  wire  dcache__EVAL_36;
  wire  dcache__EVAL_37;
  wire [63:0] dcache__EVAL_38;
  wire  dcache__EVAL_39;
  wire  dcache__EVAL_40;
  wire [2:0] dcache__EVAL_41;
  wire  dcache__EVAL_42;
  wire  dcache__EVAL_43;
  wire  dcache__EVAL_44;
  wire  dcache__EVAL_45;
  wire [7:0] dcache__EVAL_46;
  wire [5:0] dcache__EVAL_47;
  wire  dcache__EVAL_48;
  wire [1:0] dcache__EVAL_49;
  wire [31:0] dcache__EVAL_50;
  wire [1:0] dcache__EVAL_51;
  wire [31:0] dcache__EVAL_52;
  wire [1:0] dcache__EVAL_53;
  wire  dcache__EVAL_54;
  wire [31:0] dcache__EVAL_55;
  wire [1:0] dcache__EVAL_56;
  wire [2:0] dcache__EVAL_57;
  wire  dcache__EVAL_58;
  wire [63:0] dcache__EVAL_59;
  wire [31:0] dcache__EVAL_60;
  wire  dcache__EVAL_61;
  wire  dcache__EVAL_62;
  wire  dcache__EVAL_63;
  wire  dcache__EVAL_64;
  wire [3:0] dcache__EVAL_65;
  wire [2:0] dcache__EVAL_66;
  wire [29:0] dcache__EVAL_67;
  wire [31:0] dcache__EVAL_68;
  wire [31:0] dcache__EVAL_69;
  wire  dcache__EVAL_70;
  wire  dcache__EVAL_71;
  wire  dcache__EVAL_72;
  wire [31:0] dcache__EVAL_73;
  wire  dcache__EVAL_74;
  wire  dcache__EVAL_75;
  wire  dcache__EVAL_76;
  wire [3:0] dcache__EVAL_77;
  wire  dcache__EVAL_78;
  wire [31:0] dcache__EVAL_79;
  wire [3:0] dcache__EVAL_80;
  wire  dcache__EVAL_81;
  wire  dcache__EVAL_82;
  wire  dcache__EVAL_83;
  wire  dcache__EVAL_84;
  wire [1:0] dcache__EVAL_85;
  wire  dcache__EVAL_86;
  wire  dcache__EVAL_87;
  wire  dcache__EVAL_88;
  wire [1:0] dcache__EVAL_89;
  wire  dcache__EVAL_90;
  wire  dcache__EVAL_91;
  wire [63:0] dcache__EVAL_92;
  wire [1:0] dcache__EVAL_93;
  wire [31:0] dcache__EVAL_94;
  wire [29:0] dcache__EVAL_95;
  wire  dcache__EVAL_96;
  wire  dcache__EVAL_97;
  wire  dcache__EVAL_98;
  wire [3:0] dcache__EVAL_99;
  wire  dcache__EVAL_100;
  wire  dcache__EVAL_101;
  wire [29:0] dcache__EVAL_102;
  wire  dcache__EVAL_103;
  wire  dcache__EVAL_104;
  wire  dcache__EVAL_105;
  wire  dcache__EVAL_106;
  wire  dcache__EVAL_107;
  wire  dcache__EVAL_108;
  wire [31:0] dcache__EVAL_109;
  wire  dcache__EVAL_110;
  wire  dcache__EVAL_111;
  wire [1:0] dcache__EVAL_112;
  wire  dcache__EVAL_113;
  wire [1:0] dcache__EVAL_114;
  wire  dcache__EVAL_115;
  wire [31:0] dcache__EVAL_116;
  wire  dcache__EVAL_117;
  wire  dcache__EVAL_118;
  wire [4:0] dcache__EVAL_119;
  wire  dcache__EVAL_120;
  wire [31:0] dcache__EVAL_121;
  wire [31:0] dcache__EVAL_122;
  wire [2:0] dcache__EVAL_123;
  wire  dcache__EVAL_124;
  wire [31:0] dcache__EVAL_125;
  wire [2:0] dcache__EVAL_126;
  wire [31:0] dcache__EVAL_127;
  wire  dcache__EVAL_128;
  wire  dcache__EVAL_129;
  wire [31:0] dcache__EVAL_130;
  wire  dcache__EVAL_131;
  wire [1:0] dcache__EVAL_132;
  wire [5:0] dcache__EVAL_133;
  wire [2:0] dcache__EVAL_134;
  wire [4:0] dcache__EVAL_135;
  wire [31:0] dcache__EVAL_136;
  wire  dcache__EVAL_137;
  wire  dcache__EVAL_138;
  wire [31:0] dcache__EVAL_139;
  wire [1:0] dcache__EVAL_140;
  wire [1:0] dcache__EVAL_141;
  wire  dcache__EVAL_142;
  wire  dcache__EVAL_143;
  wire  dcache__EVAL_144;
  wire  dcache__EVAL_145;
  wire  dcache__EVAL_146;
  wire  dcache__EVAL_147;
  wire  dcache__EVAL_148;
  wire  dcache__EVAL_149;
  wire [29:0] dcache__EVAL_150;
  wire  intsink__EVAL;
  wire  intsink__EVAL_0;
  wire  intsink__EVAL_1;
  wire  buffer__EVAL;
  wire [3:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire [63:0] buffer__EVAL_2;
  wire [31:0] buffer__EVAL_3;
  wire [63:0] buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [3:0] buffer__EVAL_6;
  wire [2:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire [31:0] buffer__EVAL_12;
  wire [1:0] buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire [2:0] buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire  intsink_1__EVAL;
  wire  intsink_1__EVAL_0;
  wire  intsink_1__EVAL_1;
  wire  intsink_1__EVAL_2;
  wire  intsink_1__EVAL_3;
  wire  core__EVAL;
  wire  core__EVAL_0;
  wire  core__EVAL_1;
  wire [31:0] core__EVAL_2;
  wire  core__EVAL_3;
  wire  core__EVAL_4;
  wire [31:0] core__EVAL_5;
  wire [4:0] core__EVAL_6;
  wire [1:0] core__EVAL_7;
  wire  core__EVAL_8;
  wire [31:0] core__EVAL_9;
  wire [31:0] core__EVAL_10;
  wire [1:0] core__EVAL_11;
  wire  core__EVAL_12;
  wire [1:0] core__EVAL_13;
  wire [1:0] core__EVAL_14;
  wire [1:0] core__EVAL_15;
  wire  core__EVAL_16;
  wire [1:0] core__EVAL_17;
  wire [127:0] core__EVAL_18;
  wire  core__EVAL_19;
  wire  core__EVAL_20;
  wire [31:0] core__EVAL_21;
  wire  core__EVAL_22;
  wire [127:0] core__EVAL_23;
  wire  core__EVAL_24;
  wire [5:0] core__EVAL_25;
  wire  core__EVAL_26;
  wire  core__EVAL_27;
  wire  core__EVAL_28;
  wire  core__EVAL_29;
  wire  core__EVAL_30;
  wire  core__EVAL_31;
  wire  core__EVAL_32;
  wire  core__EVAL_33;
  wire  core__EVAL_34;
  wire  core__EVAL_35;
  wire  core__EVAL_36;
  wire [29:0] core__EVAL_37;
  wire [1:0] core__EVAL_38;
  wire  core__EVAL_39;
  wire  core__EVAL_40;
  wire  core__EVAL_41;
  wire  core__EVAL_42;
  wire  core__EVAL_43;
  wire [31:0] core__EVAL_44;
  wire  core__EVAL_45;
  wire [29:0] core__EVAL_46;
  wire  core__EVAL_47;
  wire  core__EVAL_48;
  wire  core__EVAL_49;
  wire  core__EVAL_50;
  wire [14:0] core__EVAL_51;
  wire  core__EVAL_52;
  wire  core__EVAL_53;
  wire  core__EVAL_54;
  wire  core__EVAL_55;
  wire  core__EVAL_56;
  wire  core__EVAL_57;
  wire  core__EVAL_58;
  wire  core__EVAL_59;
  wire  core__EVAL_60;
  wire [29:0] core__EVAL_61;
  wire [31:0] core__EVAL_62;
  wire  core__EVAL_63;
  wire [14:0] core__EVAL_64;
  wire  core__EVAL_65;
  wire [29:0] core__EVAL_66;
  wire  core__EVAL_67;
  wire [4:0] core__EVAL_68;
  wire  core__EVAL_69;
  wire  core__EVAL_70;
  wire  core__EVAL_71;
  wire  core__EVAL_72;
  wire [6:0] core__EVAL_73;
  wire  core__EVAL_74;
  wire [2:0] core__EVAL_75;
  wire  core__EVAL_76;
  wire  core__EVAL_77;
  wire  core__EVAL_78;
  wire  core__EVAL_79;
  wire  core__EVAL_80;
  wire  core__EVAL_81;
  wire  core__EVAL_82;
  wire  core__EVAL_83;
  wire [2:0] core__EVAL_84;
  wire [31:0] core__EVAL_85;
  wire  core__EVAL_86;
  wire  core__EVAL_87;
  wire [29:0] core__EVAL_88;
  wire [29:0] core__EVAL_89;
  wire  core__EVAL_90;
  wire [4:0] core__EVAL_91;
  wire  core__EVAL_92;
  wire  core__EVAL_93;
  wire [5:0] core__EVAL_94;
  wire  core__EVAL_95;
  wire [1:0] core__EVAL_96;
  wire [127:0] core__EVAL_97;
  wire  core__EVAL_98;
  wire [2:0] core__EVAL_99;
  wire  core__EVAL_100;
  wire  core__EVAL_101;
  wire  core__EVAL_102;
  wire  core__EVAL_103;
  wire  core__EVAL_104;
  wire  core__EVAL_105;
  wire  core__EVAL_106;
  wire  core__EVAL_107;
  wire  core__EVAL_108;
  wire  core__EVAL_109;
  wire [31:0] core__EVAL_110;
  wire [5:0] core__EVAL_111;
  wire  core__EVAL_112;
  wire  core__EVAL_113;
  wire  core__EVAL_114;
  wire  core__EVAL_115;
  wire  core__EVAL_116;
  wire  core__EVAL_117;
  wire  core__EVAL_118;
  wire  core__EVAL_119;
  wire  core__EVAL_120;
  wire [6:0] core__EVAL_121;
  wire  core__EVAL_122;
  wire  core__EVAL_123;
  wire  core__EVAL_124;
  wire  core__EVAL_125;
  wire [31:0] core__EVAL_126;
  wire  core__EVAL_127;
  wire  core__EVAL_128;
  wire  core__EVAL_129;
  wire  core__EVAL_130;
  wire  core__EVAL_131;
  wire [1:0] core__EVAL_132;
  wire [31:0] core__EVAL_133;
  wire  core__EVAL_134;
  wire [1:0] core__EVAL_135;
  wire  core__EVAL_136;
  wire  core__EVAL_137;
  wire [31:0] core__EVAL_138;
  wire  core__EVAL_139;
  wire  core__EVAL_140;
  wire  core__EVAL_141;
  wire  core__EVAL_142;
  wire [1:0] core__EVAL_143;
  wire  core__EVAL_144;
  wire  core__EVAL_145;
  wire  core__EVAL_146;
  wire  core__EVAL_147;
  wire  core__EVAL_148;
  wire  core__EVAL_149;
  wire  core__EVAL_150;
  wire [31:0] core__EVAL_151;
  wire  core__EVAL_152;
  wire [2:0] core__EVAL_153;
  wire [4:0] core__EVAL_154;
  wire  core__EVAL_155;
  wire  core__EVAL_156;
  wire  core__EVAL_157;
  wire [2:0] core__EVAL_158;
  wire  core__EVAL_159;
  wire  core__EVAL_160;
  wire [1:0] core__EVAL_161;
  wire [31:0] core__EVAL_162;
  wire  core__EVAL_163;
  wire  core__EVAL_164;
  wire  core__EVAL_165;
  wire [31:0] core__EVAL_166;
  wire  core__EVAL_167;
  wire  core__EVAL_168;
  wire  core__EVAL_169;
  wire  core__EVAL_170;
  wire [4:0] core__EVAL_171;
  wire  core__EVAL_172;
  wire  core__EVAL_173;
  wire  core__EVAL_174;
  wire  core__EVAL_175;
  wire  core__EVAL_176;
  wire  core__EVAL_177;
  wire [1:0] core__EVAL_178;
  wire  core__EVAL_179;
  wire [4:0] core__EVAL_180;
  wire  core__EVAL_181;
  wire  core__EVAL_182;
  wire [2:0] core__EVAL_183;
  wire  core__EVAL_184;
  wire [127:0] core__EVAL_185;
  wire  core__EVAL_186;
  wire [31:0] core__EVAL_187;
  wire  core__EVAL_188;
  wire [31:0] core__EVAL_189;
  wire  core__EVAL_190;
  wire [4:0] core__EVAL_191;
  wire  core__EVAL_192;
  wire  core__EVAL_193;
  wire [31:0] core__EVAL_194;
  wire [31:0] core__EVAL_195;
  wire  core__EVAL_196;
  wire  core__EVAL_197;
  wire  core__EVAL_198;
  wire [31:0] core__EVAL_199;
  wire [31:0] core__EVAL_200;
  wire  core__EVAL_201;
  wire [1:0] core__EVAL_202;
  wire [4:0] core__EVAL_203;
  wire  core__EVAL_204;
  wire  core__EVAL_205;
  wire  core__EVAL_206;
  wire  core__EVAL_207;
  wire [2:0] core__EVAL_208;
  wire [31:0] core__EVAL_209;
  wire  core__EVAL_210;
  wire [1:0] core__EVAL_211;
  wire  core__EVAL_212;
  wire  core__EVAL_213;
  wire  core__EVAL_214;
  wire  core__EVAL_215;
  wire  core__EVAL_216;
  wire [1:0] core__EVAL_217;
  wire  core__EVAL_218;
  wire  core__EVAL_219;
  wire  core__EVAL_220;
  wire [1:0] core__EVAL_221;
  wire [2:0] core__EVAL_222;
  wire  core__EVAL_223;
  wire  core__EVAL_224;
  wire  core__EVAL_225;
  wire  core__EVAL_226;
  wire  core__EVAL_227;
  wire  core__EVAL_228;
  wire  core__EVAL_229;
  wire [29:0] core__EVAL_230;
  wire  core__EVAL_231;
  wire  core__EVAL_232;
  wire  core__EVAL_233;
  wire [31:0] core__EVAL_234;
  wire  core__EVAL_235;
  wire  core__EVAL_236;
  wire  core__EVAL_237;
  wire [31:0] core__EVAL_238;
  wire  core__EVAL_239;
  wire [31:0] core__EVAL_240;
  wire [1:0] core__EVAL_241;
  wire  core__EVAL_242;
  wire  core__EVAL_243;
  wire  core__EVAL_244;
  wire  core__EVAL_245;
  wire  core__EVAL_246;
  wire  core__EVAL_247;
  wire [4:0] core__EVAL_248;
  wire  core__EVAL_249;
  wire  core__EVAL_250;
  wire  core__EVAL_251;
  wire  core__EVAL_252;
  wire  core__EVAL_253;
  wire  core__EVAL_254;
  wire  core__EVAL_255;
  wire [1:0] core__EVAL_256;
  wire  core__EVAL_257;
  wire  core__EVAL_258;
  wire  core__EVAL_259;
  wire  core__EVAL_260;
  wire  core__EVAL_261;
  wire [1:0] core__EVAL_262;
  wire [31:0] core__EVAL_263;
  wire [29:0] core__EVAL_264;
  wire  core__EVAL_265;
  wire [31:0] core__EVAL_266;
  wire  core__EVAL_267;
  wire  core__EVAL_268;
  wire [31:0] core__EVAL_269;
  wire [31:0] core__EVAL_270;
  wire  core__EVAL_271;
  wire  core__EVAL_272;
  wire [31:0] core__EVAL_273;
  wire [4:0] core__EVAL_274;
  wire [14:0] core__EVAL_275;
  wire  core__EVAL_276;
  wire  core__EVAL_277;
  wire  core__EVAL_278;
  wire  core__EVAL_279;
  wire [31:0] widget_1__EVAL;
  wire  widget_1__EVAL_0;
  wire [31:0] widget_1__EVAL_1;
  wire [2:0] widget_1__EVAL_2;
  wire [2:0] widget_1__EVAL_3;
  wire  widget_1__EVAL_4;
  wire [2:0] widget_1__EVAL_5;
  wire  widget_1__EVAL_6;
  wire [2:0] widget_1__EVAL_7;
  wire  widget_1__EVAL_8;
  wire [2:0] widget_1__EVAL_9;
  wire  widget_1__EVAL_10;
  wire  widget_1__EVAL_11;
  wire  widget_1__EVAL_12;
  wire [2:0] widget_1__EVAL_13;
  wire [2:0] widget_1__EVAL_14;
  wire  widget_1__EVAL_15;
  wire [63:0] widget_1__EVAL_16;
  wire  widget_1__EVAL_17;
  wire [2:0] widget_1__EVAL_18;
  wire [7:0] widget_1__EVAL_19;
  wire [2:0] widget_1__EVAL_20;
  wire [2:0] widget_1__EVAL_21;
  wire  widget_1__EVAL_22;
  wire [24:0] widget_1__EVAL_23;
  wire [63:0] widget_1__EVAL_24;
  wire [2:0] widget_1__EVAL_25;
  wire  widget_1__EVAL_26;
  wire [3:0] widget_1__EVAL_27;
  wire [2:0] widget_1__EVAL_28;
  wire [24:0] widget_1__EVAL_29;
  wire [2:0] widget_1__EVAL_30;
  wire  widget_1__EVAL_31;
  wire [2:0] widget_1__EVAL_32;
  wire [2:0] filter__EVAL;
  wire [2:0] filter__EVAL_0;
  wire  filter__EVAL_1;
  wire [7:0] filter__EVAL_2;
  wire  filter__EVAL_3;
  wire  filter__EVAL_4;
  wire [31:0] filter__EVAL_5;
  wire [2:0] filter__EVAL_6;
  wire  filter__EVAL_7;
  wire  filter__EVAL_8;
  wire  filter__EVAL_9;
  wire [3:0] filter__EVAL_10;
  wire [1:0] filter__EVAL_11;
  wire  filter__EVAL_12;
  wire [2:0] filter__EVAL_13;
  wire  filter__EVAL_14;
  wire [1:0] filter__EVAL_15;
  wire  filter__EVAL_16;
  wire  filter__EVAL_17;
  wire [31:0] filter__EVAL_18;
  wire [2:0] filter__EVAL_19;
  wire  filter__EVAL_20;
  wire  filter__EVAL_21;
  wire  filter__EVAL_22;
  wire  filter__EVAL_23;
  wire  filter__EVAL_24;
  wire [3:0] filter__EVAL_25;
  wire [1:0] filter__EVAL_26;
  wire  filter__EVAL_27;
  wire [31:0] filter__EVAL_28;
  wire [2:0] filter__EVAL_29;
  wire [63:0] filter__EVAL_30;
  wire [2:0] filter__EVAL_31;
  wire [3:0] filter__EVAL_32;
  wire [63:0] filter__EVAL_33;
  wire [2:0] filter__EVAL_34;
  wire [63:0] filter__EVAL_35;
  wire [3:0] filter__EVAL_36;
  wire [63:0] filter__EVAL_37;
  wire  filter__EVAL_38;
  wire  filter__EVAL_39;
  wire [2:0] filter__EVAL_40;
  wire [1:0] filter__EVAL_41;
  wire  filter__EVAL_42;
  wire [2:0] filter__EVAL_43;
  wire  filter__EVAL_44;
  wire  filter__EVAL_45;
  wire  filter__EVAL_46;
  wire [2:0] filter__EVAL_47;
  wire  filter__EVAL_48;
  wire  filter__EVAL_49;
  wire  filter__EVAL_50;
  wire [2:0] filter__EVAL_51;
  wire [3:0] filter__EVAL_52;
  wire  filter__EVAL_53;
  wire  filter__EVAL_54;
  wire  filter__EVAL_55;
  wire [31:0] filter__EVAL_56;
  wire  filter__EVAL_57;
  wire [2:0] filter__EVAL_58;
  wire  filter__EVAL_59;
  wire  filter__EVAL_60;
  wire [3:0] filter__EVAL_61;
  wire  filter__EVAL_62;
  wire [63:0] filter__EVAL_63;
  wire [2:0] filter__EVAL_64;
  wire [63:0] filter__EVAL_65;
  wire [31:0] filter__EVAL_66;
  wire  filter__EVAL_67;
  wire [7:0] filter__EVAL_68;
  wire [31:0] filter__EVAL_69;
  wire [2:0] filter__EVAL_70;
  wire [2:0] filter__EVAL_71;
  wire  filter__EVAL_72;
  wire  intsink_2__EVAL;
  wire  intsink_2__EVAL_0;
  wire  intsink_2__EVAL_1;
  wire  FormMicroOps__EVAL;
  wire [4:0] FormMicroOps__EVAL_0;
  wire  FormMicroOps__EVAL_1;
  wire [127:0] FormMicroOps__EVAL_2;
  wire  FormMicroOps__EVAL_3;
  wire  FormMicroOps__EVAL_4;
  wire  FormMicroOps__EVAL_5;
  wire  FormMicroOps__EVAL_6;
  wire  FormMicroOps__EVAL_7;
  wire [8:0] FormMicroOps__EVAL_8;
  wire [1:0] FormMicroOps__EVAL_9;
  wire [2:0] FormMicroOps__EVAL_10;
  wire  FormMicroOps__EVAL_11;
  wire  FormMicroOps__EVAL_12;
  wire  FormMicroOps__EVAL_13;
  wire  FormMicroOps__EVAL_14;
  wire [1:0] FormMicroOps__EVAL_15;
  wire  FormMicroOps__EVAL_16;
  wire  FormMicroOps__EVAL_17;
  wire  FormMicroOps__EVAL_18;
  wire  FormMicroOps__EVAL_19;
  wire  FormMicroOps__EVAL_20;
  wire  FormMicroOps__EVAL_21;
  wire  FormMicroOps__EVAL_22;
  wire  FormMicroOps__EVAL_23;
  wire  FormMicroOps__EVAL_24;
  wire [1:0] FormMicroOps__EVAL_25;
  wire  FormMicroOps__EVAL_26;
  wire [31:0] FormMicroOps__EVAL_27;
  wire  FormMicroOps__EVAL_28;
  wire  FormMicroOps__EVAL_29;
  wire [1:0] FormMicroOps__EVAL_30;
  wire  FormMicroOps__EVAL_31;
  wire  FormMicroOps__EVAL_32;
  wire [63:0] FormMicroOps__EVAL_33;
  wire  FormMicroOps__EVAL_34;
  wire  FormMicroOps__EVAL_35;
  wire  FormMicroOps__EVAL_36;
  wire  FormMicroOps__EVAL_37;
  wire [4:0] FormMicroOps__EVAL_38;
  wire  FormMicroOps__EVAL_39;
  wire  FormMicroOps__EVAL_40;
  wire [4:0] FormMicroOps__EVAL_41;
  wire  FormMicroOps__EVAL_42;
  wire [2:0] FormMicroOps__EVAL_43;
  wire [31:0] FormMicroOps__EVAL_44;
  wire  FormMicroOps__EVAL_45;
  wire  FormMicroOps__EVAL_46;
  wire  FormMicroOps__EVAL_47;
  wire  FormMicroOps__EVAL_48;
  wire  FormMicroOps__EVAL_49;
  wire  FormMicroOps__EVAL_50;
  wire  FormMicroOps__EVAL_51;
  wire  FormMicroOps__EVAL_52;
  wire  FormMicroOps__EVAL_53;
  wire  FormMicroOps__EVAL_54;
  wire  FormMicroOps__EVAL_55;
  wire [1:0] FormMicroOps__EVAL_56;
  wire  FormMicroOps__EVAL_57;
  wire  FormMicroOps__EVAL_58;
  wire [8:0] FormMicroOps__EVAL_59;
  wire  FormMicroOps__EVAL_60;
  wire  FormMicroOps__EVAL_61;
  wire  FormMicroOps__EVAL_62;
  wire [4:0] FormMicroOps__EVAL_63;
  wire  FormMicroOps__EVAL_64;
  wire  FormMicroOps__EVAL_65;
  wire  FormMicroOps__EVAL_66;
  wire  FormMicroOps__EVAL_67;
  wire  FormMicroOps__EVAL_68;
  wire  FormMicroOps__EVAL_69;
  wire  FormMicroOps__EVAL_70;
  wire  FormMicroOps__EVAL_71;
  wire  FormMicroOps__EVAL_72;
  wire  FormMicroOps__EVAL_73;
  wire  FormMicroOps__EVAL_74;
  wire  FormMicroOps__EVAL_75;
  wire  FormMicroOps__EVAL_76;
  wire  FormMicroOps__EVAL_77;
  wire  FormMicroOps__EVAL_78;
  wire  FormMicroOps__EVAL_79;
  wire [14:0] FormMicroOps__EVAL_80;
  wire  FormMicroOps__EVAL_81;
  wire [2:0] FormMicroOps__EVAL_82;
  wire  FormMicroOps__EVAL_83;
  wire  FormMicroOps__EVAL_84;
  wire  FormMicroOps__EVAL_85;
  wire  FormMicroOps__EVAL_86;
  wire  FormMicroOps__EVAL_87;
  wire [6:0] FormMicroOps__EVAL_88;
  wire  FormMicroOps__EVAL_89;
  wire  FormMicroOps__EVAL_90;
  wire  FormMicroOps__EVAL_91;
  wire [1:0] FormMicroOps__EVAL_92;
  wire [14:0] FormMicroOps__EVAL_93;
  wire [8:0] FormMicroOps__EVAL_94;
  wire  FormMicroOps__EVAL_95;
  wire [4:0] FormMicroOps__EVAL_96;
  wire  FormMicroOps__EVAL_97;
  wire [1:0] FormMicroOps__EVAL_98;
  wire  FormMicroOps__EVAL_99;
  wire [2:0] FormMicroOps__EVAL_100;
  wire  FormMicroOps__EVAL_101;
  wire [31:0] FormMicroOps__EVAL_102;
  wire  FormMicroOps__EVAL_103;
  wire  FormMicroOps__EVAL_104;
  wire  FormMicroOps__EVAL_105;
  wire  FormMicroOps__EVAL_106;
  wire  FormMicroOps__EVAL_107;
  wire [14:0] FormMicroOps__EVAL_108;
  wire  FormMicroOps__EVAL_109;
  wire  FormMicroOps__EVAL_110;
  wire [4:0] FormMicroOps__EVAL_111;
  wire  FormMicroOps__EVAL_112;
  wire  FormMicroOps__EVAL_113;
  wire  FormMicroOps__EVAL_114;
  wire  FormMicroOps__EVAL_115;
  wire  FormMicroOps__EVAL_116;
  wire [127:0] FormMicroOps__EVAL_117;
  wire  FormMicroOps__EVAL_118;
  wire [31:0] FormMicroOps__EVAL_119;
  wire  FormMicroOps__EVAL_120;
  wire  FormMicroOps__EVAL_121;
  wire  FormMicroOps__EVAL_122;
  wire [4:0] FormMicroOps__EVAL_123;
  wire  FormMicroOps__EVAL_124;
  wire [127:0] FormMicroOps__EVAL_125;
  wire [31:0] FormMicroOps__EVAL_126;
  wire  FormMicroOps__EVAL_127;
  wire  FormMicroOps__EVAL_128;
  wire  FormMicroOps__EVAL_129;
  wire [31:0] FormMicroOps__EVAL_130;
  wire [2:0] FormMicroOps__EVAL_131;
  wire  FormMicroOps__EVAL_132;
  wire  FormMicroOps__EVAL_133;
  wire  FormMicroOps__EVAL_134;
  wire  FormMicroOps__EVAL_135;
  wire [31:0] FormMicroOps__EVAL_136;
  wire [2:0] FormMicroOps__EVAL_137;
  wire  FormMicroOps__EVAL_138;
  wire [1:0] FormMicroOps__EVAL_139;
  wire  FormMicroOps__EVAL_140;
  wire  FormMicroOps__EVAL_141;
  wire  FormMicroOps__EVAL_142;
  wire  FormMicroOps__EVAL_143;
  wire  FormMicroOps__EVAL_144;
  wire  FormMicroOps__EVAL_145;
  wire [2:0] FormMicroOps__EVAL_146;
  wire  FormMicroOps__EVAL_147;
  wire [2:0] FormMicroOps__EVAL_148;
  wire  FormMicroOps__EVAL_149;
  wire [6:0] FormMicroOps__EVAL_150;
  wire  FormMicroOps__EVAL_151;
  wire [2:0] FormMicroOps__EVAL_152;
  wire  FormMicroOps__EVAL_153;
  wire  FormMicroOps__EVAL_154;
  wire  FormMicroOps__EVAL_155;
  wire  FormMicroOps__EVAL_156;
  wire  FormMicroOps__EVAL_157;
  wire [4:0] FormMicroOps__EVAL_158;
  wire  FormMicroOps__EVAL_159;
  wire  InstructionQueue__EVAL;
  wire  InstructionQueue__EVAL_0;
  wire [1:0] InstructionQueue__EVAL_1;
  wire  InstructionQueue__EVAL_2;
  wire [2:0] InstructionQueue__EVAL_3;
  wire  InstructionQueue__EVAL_4;
  wire  InstructionQueue__EVAL_5;
  wire  InstructionQueue__EVAL_6;
  wire  InstructionQueue__EVAL_7;
  wire  InstructionQueue__EVAL_8;
  wire [4:0] InstructionQueue__EVAL_9;
  wire  InstructionQueue__EVAL_10;
  wire  InstructionQueue__EVAL_11;
  wire  InstructionQueue__EVAL_12;
  wire [4:0] InstructionQueue__EVAL_13;
  wire  InstructionQueue__EVAL_14;
  wire  InstructionQueue__EVAL_15;
  wire  InstructionQueue__EVAL_16;
  wire  InstructionQueue__EVAL_17;
  wire [2:0] InstructionQueue__EVAL_18;
  wire  InstructionQueue__EVAL_19;
  wire  InstructionQueue__EVAL_20;
  wire  InstructionQueue__EVAL_21;
  wire  InstructionQueue__EVAL_22;
  wire [127:0] InstructionQueue__EVAL_23;
  wire [14:0] InstructionQueue__EVAL_24;
  wire  InstructionQueue__EVAL_25;
  wire  InstructionQueue__EVAL_26;
  wire [4:0] InstructionQueue__EVAL_27;
  wire  InstructionQueue__EVAL_28;
  wire [127:0] InstructionQueue__EVAL_29;
  wire [2:0] InstructionQueue__EVAL_30;
  wire [4:0] InstructionQueue__EVAL_31;
  wire  InstructionQueue__EVAL_32;
  wire  InstructionQueue__EVAL_33;
  wire  InstructionQueue__EVAL_34;
  wire  InstructionQueue__EVAL_35;
  wire  InstructionQueue__EVAL_36;
  wire  InstructionQueue__EVAL_37;
  wire  InstructionQueue__EVAL_38;
  wire [14:0] InstructionQueue__EVAL_39;
  wire  InstructionQueue__EVAL_40;
  wire [14:0] InstructionQueue__EVAL_41;
  wire  InstructionQueue__EVAL_42;
  wire  InstructionQueue__EVAL_43;
  wire  InstructionQueue__EVAL_44;
  wire  InstructionQueue__EVAL_45;
  wire  InstructionQueue__EVAL_46;
  wire [2:0] InstructionQueue__EVAL_47;
  wire [4:0] InstructionQueue__EVAL_48;
  wire  InstructionQueue__EVAL_49;
  wire  InstructionQueue__EVAL_50;
  wire  InstructionQueue__EVAL_51;
  wire  InstructionQueue__EVAL_52;
  wire  InstructionQueue__EVAL_53;
  wire  InstructionQueue__EVAL_54;
  wire  InstructionQueue__EVAL_55;
  wire  InstructionQueue__EVAL_56;
  wire  InstructionQueue__EVAL_57;
  wire [4:0] InstructionQueue__EVAL_58;
  wire  InstructionQueue__EVAL_59;
  wire  InstructionQueue__EVAL_60;
  wire  InstructionQueue__EVAL_61;
  wire [4:0] InstructionQueue__EVAL_62;
  wire [6:0] InstructionQueue__EVAL_63;
  wire  InstructionQueue__EVAL_64;
  wire  InstructionQueue__EVAL_65;
  wire  InstructionQueue__EVAL_66;
  wire  InstructionQueue__EVAL_67;
  wire  InstructionQueue__EVAL_68;
  wire [1:0] InstructionQueue__EVAL_69;
  wire  InstructionQueue__EVAL_70;
  wire  InstructionQueue__EVAL_71;
  wire [8:0] InstructionQueue__EVAL_72;
  wire  InstructionQueue__EVAL_73;
  wire [4:0] InstructionQueue__EVAL_74;
  wire  InstructionQueue__EVAL_75;
  wire  InstructionQueue__EVAL_76;
  wire [31:0] InstructionQueue__EVAL_77;
  wire  InstructionQueue__EVAL_78;
  wire  InstructionQueue__EVAL_79;
  wire  InstructionQueue__EVAL_80;
  wire  InstructionQueue__EVAL_81;
  wire [2:0] InstructionQueue__EVAL_82;
  wire  InstructionQueue__EVAL_83;
  wire  InstructionQueue__EVAL_84;
  wire  InstructionQueue__EVAL_85;
  wire  InstructionQueue__EVAL_86;
  wire  InstructionQueue__EVAL_87;
  wire [4:0] InstructionQueue__EVAL_88;
  wire  InstructionQueue__EVAL_89;
  wire  InstructionQueue__EVAL_90;
  wire [4:0] InstructionQueue__EVAL_91;
  wire [2:0] InstructionQueue__EVAL_92;
  wire  InstructionQueue__EVAL_93;
  wire  InstructionQueue__EVAL_94;
  wire  InstructionQueue__EVAL_95;
  wire  InstructionQueue__EVAL_96;
  wire  InstructionQueue__EVAL_97;
  wire [127:0] InstructionQueue__EVAL_98;
  wire  InstructionQueue__EVAL_99;
  wire  InstructionQueue__EVAL_100;
  wire [2:0] InstructionQueue__EVAL_101;
  wire [31:0] InstructionQueue__EVAL_102;
  wire [1:0] InstructionQueue__EVAL_103;
  wire  InstructionQueue__EVAL_104;
  wire  InstructionQueue__EVAL_105;
  wire  InstructionQueue__EVAL_106;
  wire [8:0] InstructionQueue__EVAL_107;
  wire  InstructionQueue__EVAL_108;
  wire [4:0] InstructionQueue__EVAL_109;
  wire  InstructionQueue__EVAL_110;
  wire  InstructionQueue__EVAL_111;
  wire  InstructionQueue__EVAL_112;
  wire  InstructionQueue__EVAL_113;
  wire  InstructionQueue__EVAL_114;
  wire  InstructionQueue__EVAL_115;
  wire  InstructionQueue__EVAL_116;
  wire [4:0] InstructionQueue__EVAL_117;
  wire  InstructionQueue__EVAL_118;
  wire  InstructionQueue__EVAL_119;
  wire  InstructionQueue__EVAL_120;
  wire  InstructionQueue__EVAL_121;
  wire  InstructionQueue__EVAL_122;
  wire  InstructionQueue__EVAL_123;
  wire  InstructionQueue__EVAL_124;
  wire [14:0] InstructionQueue__EVAL_125;
  wire [2:0] InstructionQueue__EVAL_126;
  wire [31:0] InstructionQueue__EVAL_127;
  wire [2:0] InstructionQueue__EVAL_128;
  wire [6:0] InstructionQueue__EVAL_129;
  wire  InstructionQueue__EVAL_130;
  wire  InstructionQueue__EVAL_131;
  wire  InstructionQueue__EVAL_132;
  wire [4:0] InstructionQueue__EVAL_133;
  wire  InstructionQueue__EVAL_134;
  wire  InstructionQueue__EVAL_135;
  wire  InstructionQueue__EVAL_136;
  wire  InstructionQueue__EVAL_137;
  wire  InstructionQueue__EVAL_138;
  wire  InstructionQueue__EVAL_139;
  wire  InstructionQueue__EVAL_140;
  wire [4:0] InstructionQueue__EVAL_141;
  wire  InstructionQueue__EVAL_142;
  wire  InstructionQueue__EVAL_143;
  wire  InstructionQueue__EVAL_144;
  wire [1:0] InstructionQueue__EVAL_145;
  wire [31:0] InstructionQueue__EVAL_146;
  wire  InstructionQueue__EVAL_147;
  wire [6:0] InstructionQueue__EVAL_148;
  wire [2:0] InstructionQueue__EVAL_149;
  wire  InstructionQueue__EVAL_150;
  wire  InstructionQueue__EVAL_151;
  wire [127:0] InstructionQueue__EVAL_152;
  wire  InstructionQueue__EVAL_153;
  wire [4:0] InstructionQueue__EVAL_154;
  wire  InstructionQueue__EVAL_155;
  wire  InstructionQueue__EVAL_156;
  wire  InstructionQueue__EVAL_157;
  wire  InstructionQueue__EVAL_158;
  wire  InstructionQueue__EVAL_159;
  wire  InstructionQueue__EVAL_160;
  wire  InstructionQueue__EVAL_161;
  wire  InstructionQueue__EVAL_162;
  wire [2:0] InstructionQueue__EVAL_163;
  wire  InstructionQueue__EVAL_164;
  wire  InstructionQueue__EVAL_165;
  wire  InstructionQueue__EVAL_166;
  wire  InstructionQueue__EVAL_167;
  wire  InstructionQueue__EVAL_168;
  wire [4:0] InstructionQueue__EVAL_169;
  wire  InstructionQueue__EVAL_170;
  wire [6:0] InstructionQueue__EVAL_171;
  wire  InstructionQueue__EVAL_172;
  wire  InstructionQueue__EVAL_173;
  wire  InstructionQueue__EVAL_174;
  wire  InstructionQueue__EVAL_175;
  wire  InstructionQueue__EVAL_176;
  wire  InstructionQueue__EVAL_177;
  wire  InstructionQueue__EVAL_178;
  wire  InstructionQueue__EVAL_179;
  wire  InstructionQueue__EVAL_180;
  wire  InstructionQueue__EVAL_181;
  wire  InstructionQueue__EVAL_182;
  wire [2:0] InstructionQueue__EVAL_183;
  wire  InstructionQueue__EVAL_184;
  wire  InstructionQueue__EVAL_185;
  wire [31:0] tlSlaveXbar__EVAL;
  wire [31:0] tlSlaveXbar__EVAL_0;
  wire  tlSlaveXbar__EVAL_1;
  wire [24:0] tlSlaveXbar__EVAL_2;
  wire [2:0] tlSlaveXbar__EVAL_3;
  wire [2:0] tlSlaveXbar__EVAL_4;
  wire [2:0] tlSlaveXbar__EVAL_5;
  wire [1:0] tlSlaveXbar__EVAL_6;
  wire [2:0] tlSlaveXbar__EVAL_7;
  wire  tlSlaveXbar__EVAL_8;
  wire [2:0] tlSlaveXbar__EVAL_9;
  wire  tlSlaveXbar__EVAL_10;
  wire [2:0] tlSlaveXbar__EVAL_11;
  wire  tlSlaveXbar__EVAL_12;
  wire  tlSlaveXbar__EVAL_13;
  wire [31:0] tlSlaveXbar__EVAL_14;
  wire  tlSlaveXbar__EVAL_15;
  wire [3:0] tlSlaveXbar__EVAL_16;
  wire [2:0] tlSlaveXbar__EVAL_17;
  wire  tlSlaveXbar__EVAL_18;
  wire [2:0] tlSlaveXbar__EVAL_19;
  wire [6:0] tlSlaveXbar__EVAL_20;
  wire [24:0] tlSlaveXbar__EVAL_21;
  wire [6:0] tlSlaveXbar__EVAL_22;
  wire [2:0] tlSlaveXbar__EVAL_23;
  wire  tlSlaveXbar__EVAL_24;
  wire [2:0] tlSlaveXbar__EVAL_25;
  wire  tlSlaveXbar__EVAL_26;
  wire  tlSlaveXbar__EVAL_27;
  wire [2:0] tlSlaveXbar__EVAL_28;
  wire  tlSlaveXbar__EVAL_29;
  wire [6:0] tlSlaveXbar__EVAL_30;
  wire [6:0] tlSlaveXbar__EVAL_31;
  wire [6:0] tlSlaveXbar__EVAL_32;
  wire [2:0] tlSlaveXbar__EVAL_33;
  wire  tlSlaveXbar__EVAL_34;
  wire [6:0] tlSlaveXbar__EVAL_35;
  wire [3:0] tlSlaveXbar__EVAL_36;
  wire [2:0] tlSlaveXbar__EVAL_37;
  wire  tlSlaveXbar__EVAL_38;
  wire [3:0] tlSlaveXbar__EVAL_39;
  wire [31:0] tlSlaveXbar__EVAL_40;
  wire  tlSlaveXbar__EVAL_41;
  wire  tlSlaveXbar__EVAL_42;
  wire [24:0] tlSlaveXbar__EVAL_43;
  wire  tlSlaveXbar__EVAL_44;
  wire  tlSlaveXbar__EVAL_45;
  wire  tlSlaveXbar__EVAL_46;
  wire [31:0] tlSlaveXbar__EVAL_47;
  wire  tlSlaveXbar__EVAL_48;
  wire [2:0] tlSlaveXbar__EVAL_49;
  wire [31:0] tlSlaveXbar__EVAL_50;
  wire  buffer_2__EVAL;
  wire [31:0] buffer_2__EVAL_0;
  wire  buffer_2__EVAL_1;
  wire [31:0] buffer_2__EVAL_2;
  wire  buffer_2__EVAL_3;
  wire  buffer_2__EVAL_4;
  wire [2:0] buffer_2__EVAL_5;
  wire  buffer_2__EVAL_6;
  wire [2:0] buffer_2__EVAL_7;
  wire [3:0] buffer_2__EVAL_8;
  wire [7:0] buffer_2__EVAL_9;
  wire [1:0] buffer_2__EVAL_10;
  wire [63:0] buffer_2__EVAL_11;
  wire  buffer_2__EVAL_12;
  wire [2:0] buffer_2__EVAL_13;
  wire  buffer_2__EVAL_14;
  wire [3:0] buffer_2__EVAL_15;
  wire [3:0] buffer_2__EVAL_16;
  wire [63:0] buffer_2__EVAL_17;
  wire  buffer_2__EVAL_18;
  wire  buffer_2__EVAL_19;
  wire  buffer_2__EVAL_20;
  wire  buffer_2__EVAL_21;
  wire [31:0] buffer_2__EVAL_22;
  wire [7:0] buffer_2__EVAL_23;
  wire  buffer_2__EVAL_24;
  wire [2:0] buffer_2__EVAL_25;
  wire [3:0] buffer_2__EVAL_26;
  wire  buffer_2__EVAL_27;
  wire [1:0] buffer_2__EVAL_28;
  wire [3:0] buffer_2__EVAL_29;
  wire  buffer_2__EVAL_30;
  wire [2:0] buffer_2__EVAL_31;
  wire [1:0] buffer_2__EVAL_32;
  wire  buffer_2__EVAL_33;
  wire [2:0] buffer_2__EVAL_34;
  wire [3:0] buffer_2__EVAL_35;
  wire [2:0] buffer_2__EVAL_36;
  wire  buffer_2__EVAL_37;
  wire  buffer_2__EVAL_38;
  wire  buffer_2__EVAL_39;
  wire [31:0] buffer_2__EVAL_40;
  wire [3:0] buffer_2__EVAL_41;
  wire [63:0] buffer_2__EVAL_42;
  wire [63:0] buffer_2__EVAL_43;
  wire  buffer_2__EVAL_44;
  wire [31:0] buffer_2__EVAL_45;
  wire  buffer_2__EVAL_46;
  wire  buffer_2__EVAL_47;
  wire  buffer_2__EVAL_48;
  wire [1:0] buffer_2__EVAL_49;
  wire  buffer_2__EVAL_50;
  wire  buffer_2__EVAL_51;
  wire  buffer_2__EVAL_52;
  wire  buffer_2__EVAL_53;
  wire  buffer_2__EVAL_54;
  wire  buffer_2__EVAL_55;
  wire  buffer_2__EVAL_56;
  wire [3:0] buffer_2__EVAL_57;
  wire [3:0] buffer_2__EVAL_58;
  wire [31:0] buffer_2__EVAL_59;
  wire [3:0] buffer_2__EVAL_60;
  wire [2:0] buffer_2__EVAL_61;
  wire [3:0] buffer_2__EVAL_62;
  wire  buffer_2__EVAL_63;
  wire [63:0] buffer_2__EVAL_64;
  wire  buffer_2__EVAL_65;
  wire  buffer_2__EVAL_66;
  wire [2:0] buffer_2__EVAL_67;
  wire [63:0] buffer_2__EVAL_68;
  wire [3:0] buffer_2__EVAL_69;
  wire  buffer_2__EVAL_70;
  wire [2:0] buffer_2__EVAL_71;
  wire  buffer_2__EVAL_72;
  wire  buffer_1__EVAL;
  wire [3:0] buffer_1__EVAL_0;
  wire  buffer_1__EVAL_1;
  wire [24:0] buffer_1__EVAL_2;
  wire [2:0] buffer_1__EVAL_3;
  wire [31:0] buffer_1__EVAL_4;
  wire [31:0] buffer_1__EVAL_5;
  wire [2:0] buffer_1__EVAL_6;
  wire [31:0] buffer_1__EVAL_7;
  wire  buffer_1__EVAL_8;
  wire [2:0] buffer_1__EVAL_9;
  wire [7:0] buffer_1__EVAL_10;
  wire [2:0] buffer_1__EVAL_11;
  wire [3:0] buffer_1__EVAL_12;
  wire  buffer_1__EVAL_13;
  wire  buffer_1__EVAL_14;
  wire [7:0] buffer_1__EVAL_15;
  wire  buffer_1__EVAL_16;
  wire [2:0] buffer_1__EVAL_17;
  wire  buffer_1__EVAL_18;
  wire [31:0] buffer_1__EVAL_19;
  wire [7:0] buffer_1__EVAL_20;
  wire [2:0] buffer_1__EVAL_21;
  wire [2:0] buffer_1__EVAL_22;
  wire [2:0] buffer_1__EVAL_23;
  wire  buffer_1__EVAL_24;
  wire  buffer_1__EVAL_25;
  wire  buffer_1__EVAL_26;
  wire [2:0] buffer_1__EVAL_27;
  wire  buffer_1__EVAL_28;
  wire [2:0] buffer_1__EVAL_29;
  wire  buffer_1__EVAL_30;
  wire [24:0] buffer_1__EVAL_31;
  wire [7:0] buffer_1__EVAL_32;
  wire  dcacheArb__EVAL;
  wire  dcacheArb__EVAL_0;
  wire [1:0] dcacheArb__EVAL_1;
  wire [31:0] dcacheArb__EVAL_2;
  wire  dcacheArb__EVAL_3;
  wire [31:0] dcacheArb__EVAL_4;
  wire  dcacheArb__EVAL_5;
  wire  dcacheArb__EVAL_6;
  wire  dcacheArb__EVAL_7;
  wire  dcacheArb__EVAL_8;
  wire  dcacheArb__EVAL_9;
  wire  dcacheArb__EVAL_10;
  wire [4:0] dcacheArb__EVAL_11;
  wire [31:0] dcacheArb__EVAL_12;
  wire  dcacheArb__EVAL_13;
  wire  dcacheArb__EVAL_14;
  wire  dcacheArb__EVAL_15;
  wire  dcacheArb__EVAL_16;
  wire [31:0] dcacheArb__EVAL_17;
  wire  dcacheArb__EVAL_18;
  wire [31:0] dcacheArb__EVAL_19;
  wire  dcacheArb__EVAL_20;
  wire  dcacheArb__EVAL_21;
  wire  dcacheArb__EVAL_22;
  wire [31:0] dcacheArb__EVAL_23;
  wire  dcacheArb__EVAL_24;
  wire  dcacheArb__EVAL_25;
  wire  dcacheArb__EVAL_26;
  wire  dcacheArb__EVAL_27;
  wire  dcacheArb__EVAL_28;
  wire  dcacheArb__EVAL_29;
  wire  dcacheArb__EVAL_30;
  wire  dcacheArb__EVAL_31;
  wire [31:0] dcacheArb__EVAL_32;
  wire  dcacheArb__EVAL_33;
  wire  dcacheArb__EVAL_34;
  wire [5:0] dcacheArb__EVAL_35;
  wire [31:0] dcacheArb__EVAL_36;
  wire [5:0] dcacheArb__EVAL_37;
  wire [5:0] dcacheArb__EVAL_38;
  wire  dcacheArb__EVAL_39;
  wire  dcacheArb__EVAL_40;
  wire  dcacheArb__EVAL_41;
  wire  dcacheArb__EVAL_42;
  wire  dcacheArb__EVAL_43;
  wire  dcacheArb__EVAL_44;
  wire [4:0] dcacheArb__EVAL_45;
  wire  dcacheArb__EVAL_46;
  wire  dcacheArb__EVAL_47;
  wire  dcacheArb__EVAL_48;
  wire  dcacheArb__EVAL_49;
  wire  dcacheArb__EVAL_50;
  wire  dcacheArb__EVAL_51;
  wire  dcacheArb__EVAL_52;
  wire  dcacheArb__EVAL_53;
  wire  dcacheArb__EVAL_54;
  wire  dcacheArb__EVAL_55;
  wire  dcacheArb__EVAL_56;
  wire  dcacheArb__EVAL_57;
  wire  dcacheArb__EVAL_58;
  wire  dcacheArb__EVAL_59;
  wire  dcacheArb__EVAL_60;
  wire  dcacheArb__EVAL_61;
  wire [31:0] dcacheArb__EVAL_62;
  wire  dcacheArb__EVAL_63;
  wire  dcacheArb__EVAL_64;
  wire [31:0] dcacheArb__EVAL_65;
  wire  dcacheArb__EVAL_66;
  wire  dcacheArb__EVAL_67;
  wire  dcacheArb__EVAL_68;
  wire [31:0] dcacheArb__EVAL_69;
  wire [31:0] dcacheArb__EVAL_70;
  wire [4:0] dcacheArb__EVAL_71;
  wire [1:0] dcacheArb__EVAL_72;
  wire  dcacheArb__EVAL_73;
  wire  dcacheArb__EVAL_74;
  wire  dcacheArb__EVAL_75;
  wire [5:0] dcacheArb__EVAL_76;
  wire  dcacheArb__EVAL_77;
  wire  dcacheArb__EVAL_78;
  wire [1:0] dcacheArb__EVAL_79;
  wire  dcacheArb__EVAL_80;
  wire [5:0] dcacheArb__EVAL_81;
  wire  dcacheArb__EVAL_82;
  wire [5:0] dcacheArb__EVAL_83;
  wire [4:0] dcacheArb__EVAL_84;
  wire [1:0] dcacheArb__EVAL_85;
  wire  dcacheArb__EVAL_86;
  wire  dcacheArb__EVAL_87;
  wire  dcacheArb__EVAL_88;
  wire  dcacheArb__EVAL_89;
  wire  dcacheArb__EVAL_90;
  wire  buffer_3__EVAL;
  wire [2:0] buffer_3__EVAL_0;
  wire [2:0] buffer_3__EVAL_1;
  wire [6:0] buffer_3__EVAL_2;
  wire [3:0] buffer_3__EVAL_3;
  wire [1:0] buffer_3__EVAL_4;
  wire [1:0] buffer_3__EVAL_5;
  wire [24:0] buffer_3__EVAL_6;
  wire  buffer_3__EVAL_7;
  wire  buffer_3__EVAL_8;
  wire  buffer_3__EVAL_9;
  wire [2:0] buffer_3__EVAL_10;
  wire  buffer_3__EVAL_11;
  wire  buffer_3__EVAL_12;
  wire  buffer_3__EVAL_13;
  wire [6:0] buffer_3__EVAL_14;
  wire [2:0] buffer_3__EVAL_15;
  wire [31:0] buffer_3__EVAL_16;
  wire [2:0] buffer_3__EVAL_17;
  wire [6:0] buffer_3__EVAL_18;
  wire  buffer_3__EVAL_19;
  wire  buffer_3__EVAL_20;
  wire [24:0] buffer_3__EVAL_21;
  wire  buffer_3__EVAL_22;
  wire  buffer_3__EVAL_23;
  wire [6:0] buffer_3__EVAL_24;
  wire [31:0] buffer_3__EVAL_25;
  wire  buffer_3__EVAL_26;
  wire  buffer_3__EVAL_27;
  wire  buffer_3__EVAL_28;
  wire [3:0] buffer_3__EVAL_29;
  wire [2:0] buffer_3__EVAL_30;
  wire [2:0] buffer_3__EVAL_31;
  wire [31:0] buffer_3__EVAL_32;
  wire [31:0] buffer_3__EVAL_33;
  wire [2:0] buffer_3__EVAL_34;
  wire  buffer_3__EVAL_35;
  wire [2:0] buffer_3__EVAL_36;
  wire [2:0] buffer_3__EVAL_37;
  wire  buffer_3__EVAL_38;
  wire [63:0] coreXbar__EVAL;
  wire [2:0] coreXbar__EVAL_0;
  wire [31:0] coreXbar__EVAL_1;
  wire  coreXbar__EVAL_2;
  wire [2:0] coreXbar__EVAL_3;
  wire [63:0] coreXbar__EVAL_4;
  wire  coreXbar__EVAL_5;
  wire [3:0] coreXbar__EVAL_6;
  wire  coreXbar__EVAL_7;
  wire [3:0] coreXbar__EVAL_8;
  wire [2:0] coreXbar__EVAL_9;
  wire  coreXbar__EVAL_10;
  wire [2:0] coreXbar__EVAL_11;
  wire [7:0] coreXbar__EVAL_12;
  wire  coreXbar__EVAL_13;
  wire  coreXbar__EVAL_14;
  wire  coreXbar__EVAL_15;
  wire  coreXbar__EVAL_16;
  wire [2:0] coreXbar__EVAL_17;
  wire [7:0] coreXbar__EVAL_18;
  wire  coreXbar__EVAL_19;
  wire  coreXbar__EVAL_20;
  wire  coreXbar__EVAL_21;
  wire [2:0] coreXbar__EVAL_22;
  wire  coreXbar__EVAL_23;
  wire  coreXbar__EVAL_24;
  wire [3:0] coreXbar__EVAL_25;
  wire  coreXbar__EVAL_26;
  wire  coreXbar__EVAL_27;
  wire  coreXbar__EVAL_28;
  wire [2:0] coreXbar__EVAL_29;
  wire  coreXbar__EVAL_30;
  wire [2:0] coreXbar__EVAL_31;
  wire [31:0] coreXbar__EVAL_32;
  wire [3:0] coreXbar__EVAL_33;
  wire [2:0] coreXbar__EVAL_34;
  wire [31:0] coreXbar__EVAL_35;
  wire  coreXbar__EVAL_36;
  wire [63:0] coreXbar__EVAL_37;
  wire [63:0] coreXbar__EVAL_38;
  wire  coreXbar__EVAL_39;
  wire [2:0] coreXbar__EVAL_40;
  wire  coreXbar__EVAL_41;
  wire  coreXbar__EVAL_42;
  wire [63:0] coreXbar__EVAL_43;
  wire [63:0] coreXbar__EVAL_44;
  wire  coreXbar__EVAL_45;
  wire [3:0] coreXbar__EVAL_46;
  wire  coreXbar__EVAL_47;
  wire [63:0] coreXbar__EVAL_48;
  wire [2:0] coreXbar__EVAL_49;
  wire [1:0] coreXbar__EVAL_50;
  wire  coreXbar__EVAL_51;
  wire [2:0] coreXbar__EVAL_52;
  wire  coreXbar__EVAL_53;
  wire [2:0] coreXbar__EVAL_54;
  wire [7:0] coreXbar__EVAL_55;
  wire  coreXbar__EVAL_56;
  wire [2:0] coreXbar__EVAL_57;
  wire  coreXbar__EVAL_58;
  wire  coreXbar__EVAL_59;
  wire  coreXbar__EVAL_60;
  wire [1:0] coreXbar__EVAL_61;
  wire  coreXbar__EVAL_62;
  wire [1:0] coreXbar__EVAL_63;
  wire [2:0] coreXbar__EVAL_64;
  wire [2:0] coreXbar__EVAL_65;
  wire [2:0] coreXbar__EVAL_66;
  wire  coreXbar__EVAL_67;
  wire  coreXbar__EVAL_68;
  wire [2:0] coreXbar__EVAL_69;
  wire [63:0] coreXbar__EVAL_70;
  wire [31:0] coreXbar__EVAL_71;
  wire  coreXbar__EVAL_72;
  wire [1:0] coreXbar__EVAL_73;
  wire [2:0] coreXbar__EVAL_74;
  wire  coreXbar__EVAL_75;
  wire [24:0] coreXbar__EVAL_76;
  wire  coreXbar__EVAL_77;
  wire [31:0] coreXbar__EVAL_78;
  wire  coreXbar__EVAL_79;
  wire [2:0] coreXbar__EVAL_80;
  wire [2:0] coreXbar__EVAL_81;
  wire [2:0] coreXbar__EVAL_82;
  wire [2:0] coreXbar__EVAL_83;
  wire [31:0] coreXbar__EVAL_84;
  wire [3:0] coreXbar__EVAL_85;
  wire  coreXbar__EVAL_86;
  wire  coreXbar__EVAL_87;
  wire  coreXbar__EVAL_88;
  wire  intXbar__EVAL;
  wire  intXbar__EVAL_0;
  wire  intXbar__EVAL_1;
  wire  intXbar__EVAL_2;
  wire  intXbar__EVAL_3;
  wire  intXbar__EVAL_4;
  wire  intXbar__EVAL_5;
  wire  intXbar__EVAL_6;
  wire [31:0] tlMasterXbar__EVAL;
  wire [1:0] tlMasterXbar__EVAL_0;
  wire  tlMasterXbar__EVAL_1;
  wire  tlMasterXbar__EVAL_2;
  wire [2:0] tlMasterXbar__EVAL_3;
  wire  tlMasterXbar__EVAL_4;
  wire [2:0] tlMasterXbar__EVAL_5;
  wire [63:0] tlMasterXbar__EVAL_6;
  wire [3:0] tlMasterXbar__EVAL_7;
  wire [2:0] tlMasterXbar__EVAL_8;
  wire  tlMasterXbar__EVAL_9;
  wire  tlMasterXbar__EVAL_10;
  wire [2:0] tlMasterXbar__EVAL_11;
  wire [63:0] tlMasterXbar__EVAL_12;
  wire  tlMasterXbar__EVAL_13;
  wire [3:0] tlMasterXbar__EVAL_14;
  wire [63:0] tlMasterXbar__EVAL_15;
  wire [2:0] tlMasterXbar__EVAL_16;
  wire [31:0] tlMasterXbar__EVAL_17;
  wire [2:0] tlMasterXbar__EVAL_18;
  wire  tlMasterXbar__EVAL_19;
  wire [3:0] tlMasterXbar__EVAL_20;
  wire  tlMasterXbar__EVAL_21;
  wire [31:0] tlMasterXbar__EVAL_22;
  wire  tlMasterXbar__EVAL_23;
  wire  tlMasterXbar__EVAL_24;
  wire [31:0] tlMasterXbar__EVAL_25;
  wire [3:0] tlMasterXbar__EVAL_26;
  wire  tlMasterXbar__EVAL_27;
  wire  tlMasterXbar__EVAL_28;
  wire [2:0] tlMasterXbar__EVAL_29;
  wire [3:0] tlMasterXbar__EVAL_30;
  wire [2:0] tlMasterXbar__EVAL_31;
  wire [3:0] tlMasterXbar__EVAL_32;
  wire  tlMasterXbar__EVAL_33;
  wire  tlMasterXbar__EVAL_34;
  wire [3:0] tlMasterXbar__EVAL_35;
  wire  tlMasterXbar__EVAL_36;
  wire [63:0] tlMasterXbar__EVAL_37;
  wire [1:0] tlMasterXbar__EVAL_38;
  wire  tlMasterXbar__EVAL_39;
  wire  tlMasterXbar__EVAL_40;
  wire  tlMasterXbar__EVAL_41;
  wire [63:0] tlMasterXbar__EVAL_42;
  wire  tlMasterXbar__EVAL_43;
  wire  tlMasterXbar__EVAL_44;
  wire  tlMasterXbar__EVAL_45;
  wire [3:0] tlMasterXbar__EVAL_46;
  wire  tlMasterXbar__EVAL_47;
  wire [3:0] tlMasterXbar__EVAL_48;
  wire [63:0] tlMasterXbar__EVAL_49;
  wire  tlMasterXbar__EVAL_50;
  wire  tlMasterXbar__EVAL_51;
  wire [2:0] tlMasterXbar__EVAL_52;
  wire  tlMasterXbar__EVAL_53;
  wire [3:0] tlMasterXbar__EVAL_54;
  wire  tlMasterXbar__EVAL_55;
  wire [2:0] tlMasterXbar__EVAL_56;
  wire  tlMasterXbar__EVAL_57;
  wire  tlMasterXbar__EVAL_58;
  wire  tlMasterXbar__EVAL_59;
  wire  tlMasterXbar__EVAL_60;
  wire [2:0] tlMasterXbar__EVAL_61;
  wire  tlMasterXbar__EVAL_62;
  wire [63:0] tlMasterXbar__EVAL_63;
  wire  tlMasterXbar__EVAL_64;
  wire [31:0] tlMasterXbar__EVAL_65;
  wire [7:0] tlMasterXbar__EVAL_66;
  wire  tlMasterXbar__EVAL_67;
  wire [1:0] tlMasterXbar__EVAL_68;
  wire [1:0] tlMasterXbar__EVAL_69;
  wire [31:0] tlMasterXbar__EVAL_70;
  wire  tlMasterXbar__EVAL_71;
  wire  tlMasterXbar__EVAL_72;
  wire  tlMasterXbar__EVAL_73;
  wire [2:0] tlMasterXbar__EVAL_74;
  wire  tlMasterXbar__EVAL_75;
  wire [1:0] tlMasterXbar__EVAL_76;
  wire [7:0] tlMasterXbar__EVAL_77;
  wire [2:0] tlMasterXbar__EVAL_78;
  wire [2:0] tlMasterXbar__EVAL_79;
  wire  tlMasterXbar__EVAL_80;
  wire  tlMasterXbar__EVAL_81;
  wire [31:0] tlMasterXbar__EVAL_82;
  wire  tlMasterXbar__EVAL_83;
  wire [63:0] rsource__EVAL;
  wire [31:0] rsource__EVAL_0;
  wire  rsource__EVAL_1;
  wire [2:0] rsource__EVAL_2;
  wire  rsource__EVAL_3;
  wire  rsource__EVAL_4;
  wire [3:0] rsource__EVAL_5;
  wire [63:0] rsource__EVAL_6;
  wire  rsource__EVAL_7;
  wire [3:0] rsource__EVAL_8;
  wire [1:0] rsource__EVAL_9;
  wire  rsource__EVAL_10;
  wire [3:0] rsource__EVAL_11;
  wire [3:0] rsource__EVAL_12;
  wire  rsource__EVAL_13;
  wire [63:0] rsource__EVAL_14;
  wire [63:0] rsource__EVAL_15;
  wire  rsource__EVAL_16;
  wire  rsource__EVAL_17;
  wire [1:0] rsource__EVAL_18;
  wire [31:0] rsource__EVAL_19;
  wire [3:0] rsource__EVAL_20;
  wire [3:0] rsource__EVAL_21;
  wire [3:0] rsource__EVAL_22;
  wire  rsource__EVAL_23;
  wire [1:0] rsource__EVAL_24;
  wire [3:0] rsource__EVAL_25;
  wire [3:0] rsource__EVAL_26;
  wire  rsource__EVAL_27;
  wire  rsource__EVAL_28;
  wire  rsource__EVAL_29;
  wire [63:0] rsource__EVAL_30;
  wire [7:0] rsource__EVAL_31;
  wire  rsource__EVAL_32;
  wire [31:0] rsource__EVAL_33;
  wire [3:0] rsource__EVAL_34;
  wire [63:0] rsource__EVAL_35;
  wire [2:0] rsource__EVAL_36;
  wire [2:0] rsource__EVAL_37;
  wire  rsource__EVAL_38;
  wire  rsource__EVAL_39;
  wire [7:0] rsource__EVAL_40;
  wire [1:0] rsource__EVAL_41;
  wire  rsource__EVAL_42;
  wire  rsource__EVAL_43;
  wire  rsource__EVAL_44;
  wire [1:0] rsource__EVAL_45;
  wire [2:0] rsource__EVAL_46;
  wire  rsource__EVAL_47;
  wire [3:0] rsource__EVAL_48;
  wire [31:0] rsource__EVAL_49;
  wire [1:0] rsource__EVAL_50;
  wire [1:0] rsource__EVAL_51;
  wire [1:0] rsource__EVAL_52;
  wire  rsource__EVAL_53;
  wire [2:0] rsource__EVAL_54;
  wire  rsource__EVAL_55;
  wire [2:0] rsource__EVAL_56;
  wire [1:0] rsource__EVAL_57;
  wire  rsource__EVAL_58;
  wire  rsource__EVAL_59;
  wire [63:0] rsource__EVAL_60;
  wire  rsource__EVAL_61;
  wire [31:0] rsource__EVAL_62;
  wire [3:0] rsource__EVAL_63;
  wire [3:0] rsource__EVAL_64;
  wire [1:0] rsource__EVAL_65;
  wire [1:0] rsource__EVAL_66;
  wire  rsource__EVAL_67;
  wire [31:0] rsource__EVAL_68;
  wire [2:0] rsource__EVAL_69;
  wire [1:0] rsource__EVAL_70;
  wire [31:0] rsource__EVAL_71;
  wire  rsource__EVAL_72;
  wire  rsource__EVAL_73;
  wire [2:0] rsource__EVAL_74;
  wire  rsource__EVAL_75;
  wire [63:0] rsource__EVAL_76;
  wire  rsource__EVAL_77;
  wire  rsource__EVAL_78;
  wire [31:0] rsource__EVAL_79;
  wire  rsource__EVAL_80;
  wire [2:0] rsource__EVAL_81;
  wire [2:0] rsource__EVAL_82;
  wire  rsource__EVAL_83;
  wire [2:0] rsource__EVAL_84;
  wire [3:0] rsource__EVAL_85;
  wire [1:0] rsource__EVAL_86;
  wire  rsource__EVAL_87;
  wire [3:0] rsource__EVAL_88;
  wire [63:0] rsource__EVAL_89;
  wire [3:0] rsource__EVAL_90;
  wire [2:0] rsource__EVAL_91;
  wire [3:0] rsource__EVAL_92;
  wire [1:0] rsource__EVAL_93;
  wire  rsource__EVAL_94;
  wire [31:0] rsource__EVAL_95;
  wire  rsource__EVAL_96;
  wire [2:0] rsource__EVAL_97;
  wire [2:0] rsource__EVAL_98;
  wire [1:0] rsource__EVAL_99;
  wire [7:0] rsource__EVAL_100;
  wire [1:0] rsource__EVAL_101;
  wire  rsource__EVAL_102;
  wire [2:0] rsource__EVAL_103;
  wire  rsource__EVAL_104;
  wire  rsource__EVAL_105;
  wire [3:0] rsource__EVAL_106;
  wire  rsource__EVAL_107;
  wire  rsource__EVAL_108;
  wire [2:0] fragmenter__EVAL;
  wire [63:0] fragmenter__EVAL_0;
  wire  fragmenter__EVAL_1;
  wire [6:0] fragmenter__EVAL_2;
  wire  fragmenter__EVAL_3;
  wire [11:0] fragmenter__EVAL_4;
  wire [24:0] fragmenter__EVAL_5;
  wire [7:0] fragmenter__EVAL_6;
  wire [63:0] fragmenter__EVAL_7;
  wire [2:0] fragmenter__EVAL_8;
  wire  fragmenter__EVAL_9;
  wire [7:0] fragmenter__EVAL_10;
  wire  fragmenter__EVAL_11;
  wire [2:0] fragmenter__EVAL_12;
  wire  fragmenter__EVAL_13;
  wire  fragmenter__EVAL_14;
  wire [2:0] fragmenter__EVAL_15;
  wire [6:0] fragmenter__EVAL_16;
  wire  fragmenter__EVAL_17;
  wire [1:0] fragmenter__EVAL_18;
  wire  fragmenter__EVAL_19;
  wire [11:0] fragmenter__EVAL_20;
  wire [1:0] fragmenter__EVAL_21;
  wire [2:0] fragmenter__EVAL_22;
  wire  fragmenter__EVAL_23;
  wire [63:0] fragmenter__EVAL_24;
  wire  fragmenter__EVAL_25;
  wire [2:0] fragmenter__EVAL_26;
  wire [63:0] fragmenter__EVAL_27;
  wire [24:0] fragmenter__EVAL_28;
  wire [29:0] ptw__EVAL;
  wire  ptw__EVAL_0;
  wire  ptw__EVAL_1;
  wire  ptw__EVAL_2;
  wire [1:0] ptw__EVAL_3;
  wire  ptw__EVAL_4;
  wire  ptw__EVAL_5;
  wire [31:0] ptw__EVAL_6;
  wire [29:0] ptw__EVAL_7;
  wire  ptw__EVAL_8;
  wire [1:0] ptw__EVAL_9;
  wire [29:0] ptw__EVAL_10;
  wire  ptw__EVAL_11;
  wire [31:0] ptw__EVAL_12;
  wire [29:0] ptw__EVAL_13;
  wire [1:0] ptw__EVAL_14;
  wire [31:0] ptw__EVAL_15;
  wire  ptw__EVAL_16;
  wire [29:0] ptw__EVAL_17;
  wire  ptw__EVAL_18;
  wire  ptw__EVAL_19;
  wire  ptw__EVAL_20;
  wire [31:0] ptw__EVAL_21;
  wire [31:0] ptw__EVAL_22;
  wire  ptw__EVAL_23;
  wire  ptw__EVAL_24;
  wire [1:0] ptw__EVAL_25;
  wire [31:0] ptw__EVAL_26;
  wire [31:0] ptw__EVAL_27;
  wire [31:0] ptw__EVAL_28;
  wire  ptw__EVAL_29;
  wire  ptw__EVAL_30;
  wire [1:0] ptw__EVAL_31;
  wire  ptw__EVAL_32;
  wire  ptw__EVAL_33;
  wire  ptw__EVAL_34;
  wire [29:0] ptw__EVAL_35;
  wire  ptw__EVAL_36;
  wire  ptw__EVAL_37;
  wire [1:0] ptw__EVAL_38;
  wire  ptw__EVAL_39;
  wire  ptw__EVAL_40;
  wire [29:0] ptw__EVAL_41;
  wire  ptw__EVAL_42;
  wire  ptw__EVAL_43;
  wire  ptw__EVAL_44;
  wire  ptw__EVAL_45;
  wire  ptw__EVAL_46;
  wire  ptw__EVAL_47;
  wire  ptw__EVAL_48;
  wire [1:0] ptw__EVAL_49;
  wire [29:0] ptw__EVAL_50;
  wire  ptw__EVAL_51;
  wire  ptw__EVAL_52;
  wire [1:0] ptw__EVAL_53;
  wire  ptw__EVAL_54;
  wire [29:0] ptw__EVAL_55;
  wire [1:0] ptw__EVAL_56;
  wire  ptw__EVAL_57;
  wire  ptw__EVAL_58;
  wire  ptw__EVAL_59;
  wire  ptw__EVAL_60;
  wire  ptw__EVAL_61;
  wire [1:0] ptw__EVAL_62;
  wire [1:0] ptw__EVAL_63;
  wire  ptw__EVAL_64;
  wire [1:0] ptw__EVAL_65;
  wire  ptw__EVAL_66;
  wire  ptw__EVAL_67;
  wire  ptw__EVAL_68;
  wire [31:0] ptw__EVAL_69;
  wire  ptw__EVAL_70;
  wire [1:0] ptw__EVAL_71;
  wire  ptw__EVAL_72;
  wire  ptw__EVAL_73;
  wire [29:0] ptw__EVAL_74;
  wire  ptw__EVAL_75;
  wire  ptw__EVAL_76;
  wire  ptw__EVAL_77;
  wire [31:0] ptw__EVAL_78;
  wire [1:0] ptw__EVAL_79;
  wire  ptw__EVAL_80;
  wire  ptw__EVAL_81;
  wire [31:0] ptw__EVAL_82;
  wire  ptw__EVAL_83;
  wire [29:0] ptw__EVAL_84;
  wire  ptw__EVAL_85;
  wire  ptw__EVAL_86;
  wire  ptw__EVAL_87;
  wire [1:0] ptw__EVAL_88;
  wire [29:0] ptw__EVAL_89;
  wire [1:0] ptw__EVAL_90;
  wire  ptw__EVAL_91;
  wire  ptw__EVAL_92;
  wire  ptw__EVAL_93;
  wire [31:0] ptw__EVAL_94;
  wire  ptw__EVAL_95;
  wire [31:0] ptw__EVAL_96;
  wire  ptw__EVAL_97;
  wire [29:0] ptw__EVAL_98;
  wire [1:0] ptw__EVAL_99;
  wire  ptw__EVAL_100;
  wire  ptw__EVAL_101;
  wire [29:0] ptw__EVAL_102;
  wire [1:0] ptw__EVAL_103;
  wire [31:0] ptw__EVAL_104;
  wire  ptw__EVAL_105;
  wire [31:0] ptw__EVAL_106;
  wire [1:0] ptw__EVAL_107;
  wire [31:0] ptw__EVAL_108;
  wire  ptw__EVAL_109;
  wire  ptw__EVAL_110;
  wire  ptw__EVAL_111;
  wire [29:0] ptw__EVAL_112;
  wire  ptw__EVAL_113;
  wire  ptw__EVAL_114;
  wire  ptw__EVAL_115;
  wire  ptw__EVAL_116;
  wire [31:0] ptw__EVAL_117;
  wire  ptw__EVAL_118;
  wire [1:0] ptw__EVAL_119;
  wire  ptw__EVAL_120;
  wire  ptw__EVAL_121;
  wire [29:0] ptw__EVAL_122;
  wire  ptw__EVAL_123;
  wire  ptw__EVAL_124;
  wire [1:0] ptw__EVAL_125;
  wire  ptw__EVAL_126;
  wire  ptw__EVAL_127;
  wire  ptw__EVAL_128;
  wire [31:0] ptw__EVAL_129;
  wire [29:0] ptw__EVAL_130;
  wire  ptw__EVAL_131;
  wire [1:0] ptw__EVAL_132;
  wire [31:0] ptw__EVAL_133;
  wire  ptw__EVAL_134;
  wire  ptw__EVAL_135;
  wire [29:0] ptw__EVAL_136;
  wire  ptw__EVAL_137;
  wire  ptw__EVAL_138;
  wire  ptw__EVAL_139;
  wire  ptw__EVAL_140;
  wire [31:0] ptw__EVAL_141;
  wire  ptw__EVAL_142;
  wire  ptw__EVAL_143;
  wire  ptw__EVAL_144;
  wire [31:0] ptw__EVAL_145;
  wire  ptw__EVAL_146;
  wire  ptw__EVAL_147;
  wire [1:0] ptw__EVAL_148;
  wire  ptw__EVAL_149;
  wire [29:0] ptw__EVAL_150;
  wire [1:0] ptw__EVAL_151;
  wire [1:0] ptw__EVAL_152;
  wire  ptw__EVAL_153;
  wire [31:0] ptw__EVAL_154;
  wire [31:0] ptw__EVAL_155;
  wire [29:0] ptw__EVAL_156;
  wire [1:0] ptw__EVAL_157;
  wire  ptw__EVAL_158;
  wire [31:0] ptw__EVAL_159;
  wire [29:0] ptw__EVAL_160;
  wire [1:0] ptw__EVAL_161;
  wire  ptw__EVAL_162;
  wire  ptw__EVAL_163;
  wire  ptw__EVAL_164;
  wire [1:0] ptw__EVAL_165;
  wire  ptw__EVAL_166;
  wire  ptw__EVAL_167;
  wire [31:0] ptw__EVAL_168;
  wire [31:0] ptw__EVAL_169;
  wire  ptw__EVAL_170;
  wire [29:0] ptw__EVAL_171;
  wire  ptw__EVAL_172;
  wire [29:0] ptw__EVAL_173;
  wire  ptw__EVAL_174;
  wire [29:0] ptw__EVAL_175;
  wire  ptw__EVAL_176;
  wire  ptw__EVAL_177;
  wire  ptw__EVAL_178;
  wire  ptw__EVAL_179;
  wire [31:0] frontend__EVAL;
  wire [31:0] frontend__EVAL_0;
  wire  frontend__EVAL_1;
  wire [127:0] frontend__EVAL_2;
  wire  frontend__EVAL_3;
  wire  frontend__EVAL_4;
  wire  frontend__EVAL_5;
  wire  frontend__EVAL_6;
  wire  frontend__EVAL_7;
  wire  frontend__EVAL_8;
  wire  frontend__EVAL_9;
  wire  frontend__EVAL_10;
  wire  frontend__EVAL_11;
  wire [2:0] frontend__EVAL_12;
  wire [31:0] frontend__EVAL_13;
  wire  frontend__EVAL_14;
  wire [1:0] frontend__EVAL_15;
  wire  frontend__EVAL_16;
  wire  frontend__EVAL_17;
  wire  frontend__EVAL_18;
  wire  frontend__EVAL_19;
  wire [2:0] frontend__EVAL_20;
  wire [31:0] frontend__EVAL_21;
  wire  frontend__EVAL_22;
  wire  frontend__EVAL_23;
  wire  frontend__EVAL_24;
  wire  frontend__EVAL_25;
  wire  frontend__EVAL_26;
  wire [29:0] frontend__EVAL_27;
  wire  frontend__EVAL_28;
  wire [1:0] frontend__EVAL_29;
  wire  frontend__EVAL_30;
  wire [2:0] frontend__EVAL_31;
  wire [2:0] frontend__EVAL_32;
  wire  frontend__EVAL_33;
  wire  frontend__EVAL_34;
  wire  frontend__EVAL_35;
  wire  frontend__EVAL_36;
  wire  frontend__EVAL_37;
  wire  frontend__EVAL_38;
  wire  frontend__EVAL_39;
  wire  frontend__EVAL_40;
  wire  frontend__EVAL_41;
  wire [29:0] frontend__EVAL_42;
  wire [63:0] frontend__EVAL_43;
  wire  frontend__EVAL_44;
  wire  frontend__EVAL_45;
  wire  frontend__EVAL_46;
  wire  frontend__EVAL_47;
  wire  frontend__EVAL_48;
  wire [8:0] frontend__EVAL_49;
  wire [1:0] frontend__EVAL_50;
  wire  frontend__EVAL_51;
  wire  frontend__EVAL_52;
  wire [63:0] frontend__EVAL_53;
  wire  frontend__EVAL_54;
  wire [31:0] frontend__EVAL_55;
  wire  frontend__EVAL_56;
  wire  frontend__EVAL_57;
  wire  frontend__EVAL_58;
  wire  frontend__EVAL_59;
  wire [1:0] frontend__EVAL_60;
  wire [31:0] frontend__EVAL_61;
  wire [127:0] frontend__EVAL_62;
  wire [63:0] frontend__EVAL_63;
  wire  frontend__EVAL_64;
  wire  frontend__EVAL_65;
  wire [31:0] frontend__EVAL_66;
  wire  frontend__EVAL_67;
  wire [29:0] frontend__EVAL_68;
  wire [1:0] frontend__EVAL_69;
  wire  frontend__EVAL_70;
  wire  frontend__EVAL_71;
  wire  frontend__EVAL_72;
  wire [1:0] frontend__EVAL_73;
  wire [31:0] frontend__EVAL_74;
  wire [1:0] frontend__EVAL_75;
  wire [2:0] frontend__EVAL_76;
  wire  frontend__EVAL_77;
  wire [29:0] frontend__EVAL_78;
  wire  frontend__EVAL_79;
  wire  frontend__EVAL_80;
  wire [29:0] frontend__EVAL_81;
  wire [127:0] frontend__EVAL_82;
  wire  frontend__EVAL_83;
  wire  frontend__EVAL_84;
  wire [7:0] frontend__EVAL_85;
  wire [2:0] frontend__EVAL_86;
  wire  frontend__EVAL_87;
  wire [1:0] frontend__EVAL_88;
  wire [31:0] frontend__EVAL_89;
  wire [1:0] frontend__EVAL_90;
  wire  frontend__EVAL_91;
  wire [31:0] frontend__EVAL_92;
  wire [29:0] frontend__EVAL_93;
  wire [31:0] frontend__EVAL_94;
  wire [31:0] frontend__EVAL_95;
  wire [14:0] frontend__EVAL_96;
  wire [2:0] frontend__EVAL_97;
  wire [29:0] frontend__EVAL_98;
  wire  frontend__EVAL_99;
  wire  frontend__EVAL_100;
  wire [29:0] frontend__EVAL_101;
  wire [2:0] frontend__EVAL_102;
  wire  frontend__EVAL_103;
  wire  frontend__EVAL_104;
  wire  frontend__EVAL_105;
  wire  frontend__EVAL_106;
  wire [11:0] frontend__EVAL_107;
  wire  frontend__EVAL_108;
  wire  frontend__EVAL_109;
  wire  frontend__EVAL_110;
  wire  frontend__EVAL_111;
  wire  frontend__EVAL_112;
  wire  frontend__EVAL_113;
  wire [1:0] frontend__EVAL_114;
  wire [1:0] frontend__EVAL_115;
  wire [1:0] frontend__EVAL_116;
  wire  frontend__EVAL_117;
  wire [14:0] frontend__EVAL_118;
  wire  frontend__EVAL_119;
  wire [63:0] frontend__EVAL_120;
  wire [24:0] frontend__EVAL_121;
  wire [3:0] frontend__EVAL_122;
  wire  frontend__EVAL_123;
  wire  frontend__EVAL_124;
  wire  frontend__EVAL_125;
  wire  frontend__EVAL_126;
  wire  frontend__EVAL_127;
  wire [1:0] frontend__EVAL_128;
  wire [31:0] frontend__EVAL_129;
  wire [31:0] frontend__EVAL_130;
  wire  frontend__EVAL_131;
  wire  frontend__EVAL_132;
  wire  frontend__EVAL_133;
  wire  frontend__EVAL_134;
  wire  frontend__EVAL_135;
  wire  frontend__EVAL_136;
  wire [11:0] frontend__EVAL_137;
  wire  frontend__EVAL_138;
  wire [31:0] frontend__EVAL_139;
  wire  frontend__EVAL_140;
  wire  frontend__EVAL_141;
  wire  frontend__EVAL_142;
  wire  rsink__EVAL;
  wire [31:0] rsink__EVAL_0;
  wire [31:0] rsink__EVAL_1;
  wire  rsink__EVAL_2;
  wire [6:0] rsink__EVAL_3;
  wire [31:0] rsink__EVAL_4;
  wire [2:0] rsink__EVAL_5;
  wire [6:0] rsink__EVAL_6;
  wire  rsink__EVAL_7;
  wire [31:0] rsink__EVAL_8;
  wire [24:0] rsink__EVAL_9;
  wire [1:0] rsink__EVAL_10;
  wire [2:0] rsink__EVAL_11;
  wire [2:0] rsink__EVAL_12;
  wire [1:0] rsink__EVAL_13;
  wire  rsink__EVAL_14;
  wire [2:0] rsink__EVAL_15;
  wire  rsink__EVAL_16;
  wire  rsink__EVAL_17;
  wire  rsink__EVAL_18;
  wire [2:0] rsink__EVAL_19;
  wire  rsink__EVAL_20;
  wire  rsink__EVAL_21;
  wire [24:0] rsink__EVAL_22;
  wire [2:0] rsink__EVAL_23;
  wire [2:0] rsink__EVAL_24;
  wire [31:0] rsink__EVAL_25;
  wire [24:0] rsink__EVAL_26;
  wire  rsink__EVAL_27;
  wire [6:0] rsink__EVAL_28;
  wire [2:0] rsink__EVAL_29;
  wire [2:0] rsink__EVAL_30;
  wire [3:0] rsink__EVAL_31;
  wire [1:0] rsink__EVAL_32;
  wire  rsink__EVAL_33;
  wire [1:0] rsink__EVAL_34;
  wire [6:0] rsink__EVAL_35;
  wire [1:0] rsink__EVAL_36;
  wire [1:0] rsink__EVAL_37;
  wire  rsink__EVAL_38;
  wire [2:0] rsink__EVAL_39;
  wire  rsink__EVAL_40;
  wire [3:0] rsink__EVAL_41;
  wire [6:0] rsink__EVAL_42;
  wire [3:0] rsink__EVAL_43;
  wire  rsink__EVAL_44;
  wire [31:0] rsink__EVAL_45;
  wire [2:0] rsink__EVAL_46;
  wire  rsink__EVAL_47;
  wire [1:0] rsink__EVAL_48;
  wire [2:0] rsink__EVAL_49;
  wire  rsink__EVAL_50;
  wire  rsink__EVAL_51;
  wire [2:0] rsink__EVAL_52;
  wire  rsink__EVAL_53;
  wire [2:0] rsink__EVAL_54;
  wire [6:0] rsink__EVAL_55;
  wire  rsink__EVAL_56;
  wire  rsink__EVAL_57;
  wire  rsink__EVAL_58;
  wire  rsink__EVAL_59;
  wire [2:0] rsink__EVAL_60;
  wire [2:0] dlsXbar__EVAL;
  wire  dlsXbar__EVAL_0;
  wire [2:0] dlsXbar__EVAL_1;
  wire [31:0] dlsXbar__EVAL_2;
  wire [6:0] dlsXbar__EVAL_3;
  wire [2:0] dlsXbar__EVAL_4;
  wire  dlsXbar__EVAL_5;
  wire [2:0] dlsXbar__EVAL_6;
  wire  dlsXbar__EVAL_7;
  wire [2:0] dlsXbar__EVAL_8;
  wire  dlsXbar__EVAL_9;
  wire  dlsXbar__EVAL_10;
  wire [2:0] dlsXbar__EVAL_11;
  wire  dlsXbar__EVAL_12;
  wire [2:0] dlsXbar__EVAL_13;
  wire [31:0] dlsXbar__EVAL_14;
  wire [2:0] dlsXbar__EVAL_15;
  wire  dlsXbar__EVAL_16;
  wire  dlsXbar__EVAL_17;
  wire [31:0] dlsXbar__EVAL_18;
  wire [24:0] dlsXbar__EVAL_19;
  wire [24:0] dlsXbar__EVAL_20;
  wire [3:0] dlsXbar__EVAL_21;
  wire  dlsXbar__EVAL_22;
  wire [31:0] dlsXbar__EVAL_23;
  wire  dlsXbar__EVAL_24;
  wire [2:0] dlsXbar__EVAL_25;
  wire [3:0] dlsXbar__EVAL_26;
  wire [24:0] dlsXbar__EVAL_27;
  wire [3:0] dlsXbar__EVAL_28;
  wire [7:0] dlsXbar__EVAL_29;
  wire [2:0] dlsXbar__EVAL_30;
  wire  dlsXbar__EVAL_31;
  wire  dlsXbar__EVAL_32;
  wire  dlsXbar__EVAL_33;
  wire  dlsXbar__EVAL_34;
  wire  dlsXbar__EVAL_35;
  wire [2:0] dlsXbar__EVAL_36;
  wire [2:0] dlsXbar__EVAL_37;
  wire [2:0] dlsXbar__EVAL_38;
  wire [2:0] dlsXbar__EVAL_39;
  wire [7:0] dlsXbar__EVAL_40;
  wire [2:0] dlsXbar__EVAL_41;
  wire [31:0] dlsXbar__EVAL_42;
  wire  dlsXbar__EVAL_43;
  wire [2:0] dlsXbar__EVAL_44;
  wire [31:0] dlsXbar__EVAL_45;
  wire [6:0] dlsXbar__EVAL_46;
  wire  dlsXbar__EVAL_47;
  wire [2:0] dlsXbar__EVAL_48;
  SiFive__EVAL_249 fragmenter_1 (
    ._EVAL(fragmenter_1__EVAL),
    ._EVAL_0(fragmenter_1__EVAL_0),
    ._EVAL_1(fragmenter_1__EVAL_1),
    ._EVAL_2(fragmenter_1__EVAL_2),
    ._EVAL_3(fragmenter_1__EVAL_3),
    ._EVAL_4(fragmenter_1__EVAL_4),
    ._EVAL_5(fragmenter_1__EVAL_5),
    ._EVAL_6(fragmenter_1__EVAL_6),
    ._EVAL_7(fragmenter_1__EVAL_7),
    ._EVAL_8(fragmenter_1__EVAL_8),
    ._EVAL_9(fragmenter_1__EVAL_9),
    ._EVAL_10(fragmenter_1__EVAL_10),
    ._EVAL_11(fragmenter_1__EVAL_11),
    ._EVAL_12(fragmenter_1__EVAL_12),
    ._EVAL_13(fragmenter_1__EVAL_13),
    ._EVAL_14(fragmenter_1__EVAL_14),
    ._EVAL_15(fragmenter_1__EVAL_15),
    ._EVAL_16(fragmenter_1__EVAL_16),
    ._EVAL_17(fragmenter_1__EVAL_17),
    ._EVAL_18(fragmenter_1__EVAL_18),
    ._EVAL_19(fragmenter_1__EVAL_19),
    ._EVAL_20(fragmenter_1__EVAL_20),
    ._EVAL_21(fragmenter_1__EVAL_21),
    ._EVAL_22(fragmenter_1__EVAL_22),
    ._EVAL_23(fragmenter_1__EVAL_23),
    ._EVAL_24(fragmenter_1__EVAL_24),
    ._EVAL_25(fragmenter_1__EVAL_25),
    ._EVAL_26(fragmenter_1__EVAL_26),
    ._EVAL_27(fragmenter_1__EVAL_27),
    ._EVAL_28(fragmenter_1__EVAL_28),
    ._EVAL_29(fragmenter_1__EVAL_29),
    ._EVAL_30(fragmenter_1__EVAL_30),
    ._EVAL_31(fragmenter_1__EVAL_31),
    ._EVAL_32(fragmenter_1__EVAL_32)
  );
  SiFive__EVAL_243 dls (
    ._EVAL(dls__EVAL),
    ._EVAL_0(dls__EVAL_0),
    ._EVAL_1(dls__EVAL_1),
    ._EVAL_2(dls__EVAL_2),
    ._EVAL_3(dls__EVAL_3),
    ._EVAL_4(dls__EVAL_4),
    ._EVAL_5(dls__EVAL_5),
    ._EVAL_6(dls__EVAL_6),
    ._EVAL_7(dls__EVAL_7),
    ._EVAL_8(dls__EVAL_8),
    ._EVAL_9(dls__EVAL_9),
    ._EVAL_10(dls__EVAL_10),
    ._EVAL_11(dls__EVAL_11),
    ._EVAL_12(dls__EVAL_12),
    ._EVAL_13(dls__EVAL_13),
    ._EVAL_14(dls__EVAL_14),
    ._EVAL_15(dls__EVAL_15),
    ._EVAL_16(dls__EVAL_16)
  );
  SiFive__EVAL_238 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28)
  );
  SiFive__EVAL_259 dcache (
    ._EVAL(dcache__EVAL),
    ._EVAL_0(dcache__EVAL_0),
    ._EVAL_1(dcache__EVAL_1),
    ._EVAL_2(dcache__EVAL_2),
    ._EVAL_3(dcache__EVAL_3),
    ._EVAL_4(dcache__EVAL_4),
    ._EVAL_5(dcache__EVAL_5),
    ._EVAL_6(dcache__EVAL_6),
    ._EVAL_7(dcache__EVAL_7),
    ._EVAL_8(dcache__EVAL_8),
    ._EVAL_9(dcache__EVAL_9),
    ._EVAL_10(dcache__EVAL_10),
    ._EVAL_11(dcache__EVAL_11),
    ._EVAL_12(dcache__EVAL_12),
    ._EVAL_13(dcache__EVAL_13),
    ._EVAL_14(dcache__EVAL_14),
    ._EVAL_15(dcache__EVAL_15),
    ._EVAL_16(dcache__EVAL_16),
    ._EVAL_17(dcache__EVAL_17),
    ._EVAL_18(dcache__EVAL_18),
    ._EVAL_19(dcache__EVAL_19),
    ._EVAL_20(dcache__EVAL_20),
    ._EVAL_21(dcache__EVAL_21),
    ._EVAL_22(dcache__EVAL_22),
    ._EVAL_23(dcache__EVAL_23),
    ._EVAL_24(dcache__EVAL_24),
    ._EVAL_25(dcache__EVAL_25),
    ._EVAL_26(dcache__EVAL_26),
    ._EVAL_27(dcache__EVAL_27),
    ._EVAL_28(dcache__EVAL_28),
    ._EVAL_29(dcache__EVAL_29),
    ._EVAL_30(dcache__EVAL_30),
    ._EVAL_31(dcache__EVAL_31),
    ._EVAL_32(dcache__EVAL_32),
    ._EVAL_33(dcache__EVAL_33),
    ._EVAL_34(dcache__EVAL_34),
    ._EVAL_35(dcache__EVAL_35),
    ._EVAL_36(dcache__EVAL_36),
    ._EVAL_37(dcache__EVAL_37),
    ._EVAL_38(dcache__EVAL_38),
    ._EVAL_39(dcache__EVAL_39),
    ._EVAL_40(dcache__EVAL_40),
    ._EVAL_41(dcache__EVAL_41),
    ._EVAL_42(dcache__EVAL_42),
    ._EVAL_43(dcache__EVAL_43),
    ._EVAL_44(dcache__EVAL_44),
    ._EVAL_45(dcache__EVAL_45),
    ._EVAL_46(dcache__EVAL_46),
    ._EVAL_47(dcache__EVAL_47),
    ._EVAL_48(dcache__EVAL_48),
    ._EVAL_49(dcache__EVAL_49),
    ._EVAL_50(dcache__EVAL_50),
    ._EVAL_51(dcache__EVAL_51),
    ._EVAL_52(dcache__EVAL_52),
    ._EVAL_53(dcache__EVAL_53),
    ._EVAL_54(dcache__EVAL_54),
    ._EVAL_55(dcache__EVAL_55),
    ._EVAL_56(dcache__EVAL_56),
    ._EVAL_57(dcache__EVAL_57),
    ._EVAL_58(dcache__EVAL_58),
    ._EVAL_59(dcache__EVAL_59),
    ._EVAL_60(dcache__EVAL_60),
    ._EVAL_61(dcache__EVAL_61),
    ._EVAL_62(dcache__EVAL_62),
    ._EVAL_63(dcache__EVAL_63),
    ._EVAL_64(dcache__EVAL_64),
    ._EVAL_65(dcache__EVAL_65),
    ._EVAL_66(dcache__EVAL_66),
    ._EVAL_67(dcache__EVAL_67),
    ._EVAL_68(dcache__EVAL_68),
    ._EVAL_69(dcache__EVAL_69),
    ._EVAL_70(dcache__EVAL_70),
    ._EVAL_71(dcache__EVAL_71),
    ._EVAL_72(dcache__EVAL_72),
    ._EVAL_73(dcache__EVAL_73),
    ._EVAL_74(dcache__EVAL_74),
    ._EVAL_75(dcache__EVAL_75),
    ._EVAL_76(dcache__EVAL_76),
    ._EVAL_77(dcache__EVAL_77),
    ._EVAL_78(dcache__EVAL_78),
    ._EVAL_79(dcache__EVAL_79),
    ._EVAL_80(dcache__EVAL_80),
    ._EVAL_81(dcache__EVAL_81),
    ._EVAL_82(dcache__EVAL_82),
    ._EVAL_83(dcache__EVAL_83),
    ._EVAL_84(dcache__EVAL_84),
    ._EVAL_85(dcache__EVAL_85),
    ._EVAL_86(dcache__EVAL_86),
    ._EVAL_87(dcache__EVAL_87),
    ._EVAL_88(dcache__EVAL_88),
    ._EVAL_89(dcache__EVAL_89),
    ._EVAL_90(dcache__EVAL_90),
    ._EVAL_91(dcache__EVAL_91),
    ._EVAL_92(dcache__EVAL_92),
    ._EVAL_93(dcache__EVAL_93),
    ._EVAL_94(dcache__EVAL_94),
    ._EVAL_95(dcache__EVAL_95),
    ._EVAL_96(dcache__EVAL_96),
    ._EVAL_97(dcache__EVAL_97),
    ._EVAL_98(dcache__EVAL_98),
    ._EVAL_99(dcache__EVAL_99),
    ._EVAL_100(dcache__EVAL_100),
    ._EVAL_101(dcache__EVAL_101),
    ._EVAL_102(dcache__EVAL_102),
    ._EVAL_103(dcache__EVAL_103),
    ._EVAL_104(dcache__EVAL_104),
    ._EVAL_105(dcache__EVAL_105),
    ._EVAL_106(dcache__EVAL_106),
    ._EVAL_107(dcache__EVAL_107),
    ._EVAL_108(dcache__EVAL_108),
    ._EVAL_109(dcache__EVAL_109),
    ._EVAL_110(dcache__EVAL_110),
    ._EVAL_111(dcache__EVAL_111),
    ._EVAL_112(dcache__EVAL_112),
    ._EVAL_113(dcache__EVAL_113),
    ._EVAL_114(dcache__EVAL_114),
    ._EVAL_115(dcache__EVAL_115),
    ._EVAL_116(dcache__EVAL_116),
    ._EVAL_117(dcache__EVAL_117),
    ._EVAL_118(dcache__EVAL_118),
    ._EVAL_119(dcache__EVAL_119),
    ._EVAL_120(dcache__EVAL_120),
    ._EVAL_121(dcache__EVAL_121),
    ._EVAL_122(dcache__EVAL_122),
    ._EVAL_123(dcache__EVAL_123),
    ._EVAL_124(dcache__EVAL_124),
    ._EVAL_125(dcache__EVAL_125),
    ._EVAL_126(dcache__EVAL_126),
    ._EVAL_127(dcache__EVAL_127),
    ._EVAL_128(dcache__EVAL_128),
    ._EVAL_129(dcache__EVAL_129),
    ._EVAL_130(dcache__EVAL_130),
    ._EVAL_131(dcache__EVAL_131),
    ._EVAL_132(dcache__EVAL_132),
    ._EVAL_133(dcache__EVAL_133),
    ._EVAL_134(dcache__EVAL_134),
    ._EVAL_135(dcache__EVAL_135),
    ._EVAL_136(dcache__EVAL_136),
    ._EVAL_137(dcache__EVAL_137),
    ._EVAL_138(dcache__EVAL_138),
    ._EVAL_139(dcache__EVAL_139),
    ._EVAL_140(dcache__EVAL_140),
    ._EVAL_141(dcache__EVAL_141),
    ._EVAL_142(dcache__EVAL_142),
    ._EVAL_143(dcache__EVAL_143),
    ._EVAL_144(dcache__EVAL_144),
    ._EVAL_145(dcache__EVAL_145),
    ._EVAL_146(dcache__EVAL_146),
    ._EVAL_147(dcache__EVAL_147),
    ._EVAL_148(dcache__EVAL_148),
    ._EVAL_149(dcache__EVAL_149),
    ._EVAL_150(dcache__EVAL_150)
  );
  SiFive__EVAL_279 intsink (
    ._EVAL(intsink__EVAL),
    ._EVAL_0(intsink__EVAL_0),
    ._EVAL_1(intsink__EVAL_1)
  );
  SiFive__EVAL_240 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19)
  );
  SiFive__EVAL_281 intsink_1 (
    ._EVAL(intsink_1__EVAL),
    ._EVAL_0(intsink_1__EVAL_0),
    ._EVAL_1(intsink_1__EVAL_1),
    ._EVAL_2(intsink_1__EVAL_2),
    ._EVAL_3(intsink_1__EVAL_3)
  );
  SiFive__EVAL_307 core (
    ._EVAL(core__EVAL),
    ._EVAL_0(core__EVAL_0),
    ._EVAL_1(core__EVAL_1),
    ._EVAL_2(core__EVAL_2),
    ._EVAL_3(core__EVAL_3),
    ._EVAL_4(core__EVAL_4),
    ._EVAL_5(core__EVAL_5),
    ._EVAL_6(core__EVAL_6),
    ._EVAL_7(core__EVAL_7),
    ._EVAL_8(core__EVAL_8),
    ._EVAL_9(core__EVAL_9),
    ._EVAL_10(core__EVAL_10),
    ._EVAL_11(core__EVAL_11),
    ._EVAL_12(core__EVAL_12),
    ._EVAL_13(core__EVAL_13),
    ._EVAL_14(core__EVAL_14),
    ._EVAL_15(core__EVAL_15),
    ._EVAL_16(core__EVAL_16),
    ._EVAL_17(core__EVAL_17),
    ._EVAL_18(core__EVAL_18),
    ._EVAL_19(core__EVAL_19),
    ._EVAL_20(core__EVAL_20),
    ._EVAL_21(core__EVAL_21),
    ._EVAL_22(core__EVAL_22),
    ._EVAL_23(core__EVAL_23),
    ._EVAL_24(core__EVAL_24),
    ._EVAL_25(core__EVAL_25),
    ._EVAL_26(core__EVAL_26),
    ._EVAL_27(core__EVAL_27),
    ._EVAL_28(core__EVAL_28),
    ._EVAL_29(core__EVAL_29),
    ._EVAL_30(core__EVAL_30),
    ._EVAL_31(core__EVAL_31),
    ._EVAL_32(core__EVAL_32),
    ._EVAL_33(core__EVAL_33),
    ._EVAL_34(core__EVAL_34),
    ._EVAL_35(core__EVAL_35),
    ._EVAL_36(core__EVAL_36),
    ._EVAL_37(core__EVAL_37),
    ._EVAL_38(core__EVAL_38),
    ._EVAL_39(core__EVAL_39),
    ._EVAL_40(core__EVAL_40),
    ._EVAL_41(core__EVAL_41),
    ._EVAL_42(core__EVAL_42),
    ._EVAL_43(core__EVAL_43),
    ._EVAL_44(core__EVAL_44),
    ._EVAL_45(core__EVAL_45),
    ._EVAL_46(core__EVAL_46),
    ._EVAL_47(core__EVAL_47),
    ._EVAL_48(core__EVAL_48),
    ._EVAL_49(core__EVAL_49),
    ._EVAL_50(core__EVAL_50),
    ._EVAL_51(core__EVAL_51),
    ._EVAL_52(core__EVAL_52),
    ._EVAL_53(core__EVAL_53),
    ._EVAL_54(core__EVAL_54),
    ._EVAL_55(core__EVAL_55),
    ._EVAL_56(core__EVAL_56),
    ._EVAL_57(core__EVAL_57),
    ._EVAL_58(core__EVAL_58),
    ._EVAL_59(core__EVAL_59),
    ._EVAL_60(core__EVAL_60),
    ._EVAL_61(core__EVAL_61),
    ._EVAL_62(core__EVAL_62),
    ._EVAL_63(core__EVAL_63),
    ._EVAL_64(core__EVAL_64),
    ._EVAL_65(core__EVAL_65),
    ._EVAL_66(core__EVAL_66),
    ._EVAL_67(core__EVAL_67),
    ._EVAL_68(core__EVAL_68),
    ._EVAL_69(core__EVAL_69),
    ._EVAL_70(core__EVAL_70),
    ._EVAL_71(core__EVAL_71),
    ._EVAL_72(core__EVAL_72),
    ._EVAL_73(core__EVAL_73),
    ._EVAL_74(core__EVAL_74),
    ._EVAL_75(core__EVAL_75),
    ._EVAL_76(core__EVAL_76),
    ._EVAL_77(core__EVAL_77),
    ._EVAL_78(core__EVAL_78),
    ._EVAL_79(core__EVAL_79),
    ._EVAL_80(core__EVAL_80),
    ._EVAL_81(core__EVAL_81),
    ._EVAL_82(core__EVAL_82),
    ._EVAL_83(core__EVAL_83),
    ._EVAL_84(core__EVAL_84),
    ._EVAL_85(core__EVAL_85),
    ._EVAL_86(core__EVAL_86),
    ._EVAL_87(core__EVAL_87),
    ._EVAL_88(core__EVAL_88),
    ._EVAL_89(core__EVAL_89),
    ._EVAL_90(core__EVAL_90),
    ._EVAL_91(core__EVAL_91),
    ._EVAL_92(core__EVAL_92),
    ._EVAL_93(core__EVAL_93),
    ._EVAL_94(core__EVAL_94),
    ._EVAL_95(core__EVAL_95),
    ._EVAL_96(core__EVAL_96),
    ._EVAL_97(core__EVAL_97),
    ._EVAL_98(core__EVAL_98),
    ._EVAL_99(core__EVAL_99),
    ._EVAL_100(core__EVAL_100),
    ._EVAL_101(core__EVAL_101),
    ._EVAL_102(core__EVAL_102),
    ._EVAL_103(core__EVAL_103),
    ._EVAL_104(core__EVAL_104),
    ._EVAL_105(core__EVAL_105),
    ._EVAL_106(core__EVAL_106),
    ._EVAL_107(core__EVAL_107),
    ._EVAL_108(core__EVAL_108),
    ._EVAL_109(core__EVAL_109),
    ._EVAL_110(core__EVAL_110),
    ._EVAL_111(core__EVAL_111),
    ._EVAL_112(core__EVAL_112),
    ._EVAL_113(core__EVAL_113),
    ._EVAL_114(core__EVAL_114),
    ._EVAL_115(core__EVAL_115),
    ._EVAL_116(core__EVAL_116),
    ._EVAL_117(core__EVAL_117),
    ._EVAL_118(core__EVAL_118),
    ._EVAL_119(core__EVAL_119),
    ._EVAL_120(core__EVAL_120),
    ._EVAL_121(core__EVAL_121),
    ._EVAL_122(core__EVAL_122),
    ._EVAL_123(core__EVAL_123),
    ._EVAL_124(core__EVAL_124),
    ._EVAL_125(core__EVAL_125),
    ._EVAL_126(core__EVAL_126),
    ._EVAL_127(core__EVAL_127),
    ._EVAL_128(core__EVAL_128),
    ._EVAL_129(core__EVAL_129),
    ._EVAL_130(core__EVAL_130),
    ._EVAL_131(core__EVAL_131),
    ._EVAL_132(core__EVAL_132),
    ._EVAL_133(core__EVAL_133),
    ._EVAL_134(core__EVAL_134),
    ._EVAL_135(core__EVAL_135),
    ._EVAL_136(core__EVAL_136),
    ._EVAL_137(core__EVAL_137),
    ._EVAL_138(core__EVAL_138),
    ._EVAL_139(core__EVAL_139),
    ._EVAL_140(core__EVAL_140),
    ._EVAL_141(core__EVAL_141),
    ._EVAL_142(core__EVAL_142),
    ._EVAL_143(core__EVAL_143),
    ._EVAL_144(core__EVAL_144),
    ._EVAL_145(core__EVAL_145),
    ._EVAL_146(core__EVAL_146),
    ._EVAL_147(core__EVAL_147),
    ._EVAL_148(core__EVAL_148),
    ._EVAL_149(core__EVAL_149),
    ._EVAL_150(core__EVAL_150),
    ._EVAL_151(core__EVAL_151),
    ._EVAL_152(core__EVAL_152),
    ._EVAL_153(core__EVAL_153),
    ._EVAL_154(core__EVAL_154),
    ._EVAL_155(core__EVAL_155),
    ._EVAL_156(core__EVAL_156),
    ._EVAL_157(core__EVAL_157),
    ._EVAL_158(core__EVAL_158),
    ._EVAL_159(core__EVAL_159),
    ._EVAL_160(core__EVAL_160),
    ._EVAL_161(core__EVAL_161),
    ._EVAL_162(core__EVAL_162),
    ._EVAL_163(core__EVAL_163),
    ._EVAL_164(core__EVAL_164),
    ._EVAL_165(core__EVAL_165),
    ._EVAL_166(core__EVAL_166),
    ._EVAL_167(core__EVAL_167),
    ._EVAL_168(core__EVAL_168),
    ._EVAL_169(core__EVAL_169),
    ._EVAL_170(core__EVAL_170),
    ._EVAL_171(core__EVAL_171),
    ._EVAL_172(core__EVAL_172),
    ._EVAL_173(core__EVAL_173),
    ._EVAL_174(core__EVAL_174),
    ._EVAL_175(core__EVAL_175),
    ._EVAL_176(core__EVAL_176),
    ._EVAL_177(core__EVAL_177),
    ._EVAL_178(core__EVAL_178),
    ._EVAL_179(core__EVAL_179),
    ._EVAL_180(core__EVAL_180),
    ._EVAL_181(core__EVAL_181),
    ._EVAL_182(core__EVAL_182),
    ._EVAL_183(core__EVAL_183),
    ._EVAL_184(core__EVAL_184),
    ._EVAL_185(core__EVAL_185),
    ._EVAL_186(core__EVAL_186),
    ._EVAL_187(core__EVAL_187),
    ._EVAL_188(core__EVAL_188),
    ._EVAL_189(core__EVAL_189),
    ._EVAL_190(core__EVAL_190),
    ._EVAL_191(core__EVAL_191),
    ._EVAL_192(core__EVAL_192),
    ._EVAL_193(core__EVAL_193),
    ._EVAL_194(core__EVAL_194),
    ._EVAL_195(core__EVAL_195),
    ._EVAL_196(core__EVAL_196),
    ._EVAL_197(core__EVAL_197),
    ._EVAL_198(core__EVAL_198),
    ._EVAL_199(core__EVAL_199),
    ._EVAL_200(core__EVAL_200),
    ._EVAL_201(core__EVAL_201),
    ._EVAL_202(core__EVAL_202),
    ._EVAL_203(core__EVAL_203),
    ._EVAL_204(core__EVAL_204),
    ._EVAL_205(core__EVAL_205),
    ._EVAL_206(core__EVAL_206),
    ._EVAL_207(core__EVAL_207),
    ._EVAL_208(core__EVAL_208),
    ._EVAL_209(core__EVAL_209),
    ._EVAL_210(core__EVAL_210),
    ._EVAL_211(core__EVAL_211),
    ._EVAL_212(core__EVAL_212),
    ._EVAL_213(core__EVAL_213),
    ._EVAL_214(core__EVAL_214),
    ._EVAL_215(core__EVAL_215),
    ._EVAL_216(core__EVAL_216),
    ._EVAL_217(core__EVAL_217),
    ._EVAL_218(core__EVAL_218),
    ._EVAL_219(core__EVAL_219),
    ._EVAL_220(core__EVAL_220),
    ._EVAL_221(core__EVAL_221),
    ._EVAL_222(core__EVAL_222),
    ._EVAL_223(core__EVAL_223),
    ._EVAL_224(core__EVAL_224),
    ._EVAL_225(core__EVAL_225),
    ._EVAL_226(core__EVAL_226),
    ._EVAL_227(core__EVAL_227),
    ._EVAL_228(core__EVAL_228),
    ._EVAL_229(core__EVAL_229),
    ._EVAL_230(core__EVAL_230),
    ._EVAL_231(core__EVAL_231),
    ._EVAL_232(core__EVAL_232),
    ._EVAL_233(core__EVAL_233),
    ._EVAL_234(core__EVAL_234),
    ._EVAL_235(core__EVAL_235),
    ._EVAL_236(core__EVAL_236),
    ._EVAL_237(core__EVAL_237),
    ._EVAL_238(core__EVAL_238),
    ._EVAL_239(core__EVAL_239),
    ._EVAL_240(core__EVAL_240),
    ._EVAL_241(core__EVAL_241),
    ._EVAL_242(core__EVAL_242),
    ._EVAL_243(core__EVAL_243),
    ._EVAL_244(core__EVAL_244),
    ._EVAL_245(core__EVAL_245),
    ._EVAL_246(core__EVAL_246),
    ._EVAL_247(core__EVAL_247),
    ._EVAL_248(core__EVAL_248),
    ._EVAL_249(core__EVAL_249),
    ._EVAL_250(core__EVAL_250),
    ._EVAL_251(core__EVAL_251),
    ._EVAL_252(core__EVAL_252),
    ._EVAL_253(core__EVAL_253),
    ._EVAL_254(core__EVAL_254),
    ._EVAL_255(core__EVAL_255),
    ._EVAL_256(core__EVAL_256),
    ._EVAL_257(core__EVAL_257),
    ._EVAL_258(core__EVAL_258),
    ._EVAL_259(core__EVAL_259),
    ._EVAL_260(core__EVAL_260),
    ._EVAL_261(core__EVAL_261),
    ._EVAL_262(core__EVAL_262),
    ._EVAL_263(core__EVAL_263),
    ._EVAL_264(core__EVAL_264),
    ._EVAL_265(core__EVAL_265),
    ._EVAL_266(core__EVAL_266),
    ._EVAL_267(core__EVAL_267),
    ._EVAL_268(core__EVAL_268),
    ._EVAL_269(core__EVAL_269),
    ._EVAL_270(core__EVAL_270),
    ._EVAL_271(core__EVAL_271),
    ._EVAL_272(core__EVAL_272),
    ._EVAL_273(core__EVAL_273),
    ._EVAL_274(core__EVAL_274),
    ._EVAL_275(core__EVAL_275),
    ._EVAL_276(core__EVAL_276),
    ._EVAL_277(core__EVAL_277),
    ._EVAL_278(core__EVAL_278),
    ._EVAL_279(core__EVAL_279)
  );
  SiFive__EVAL_262 widget_1 (
    ._EVAL(widget_1__EVAL),
    ._EVAL_0(widget_1__EVAL_0),
    ._EVAL_1(widget_1__EVAL_1),
    ._EVAL_2(widget_1__EVAL_2),
    ._EVAL_3(widget_1__EVAL_3),
    ._EVAL_4(widget_1__EVAL_4),
    ._EVAL_5(widget_1__EVAL_5),
    ._EVAL_6(widget_1__EVAL_6),
    ._EVAL_7(widget_1__EVAL_7),
    ._EVAL_8(widget_1__EVAL_8),
    ._EVAL_9(widget_1__EVAL_9),
    ._EVAL_10(widget_1__EVAL_10),
    ._EVAL_11(widget_1__EVAL_11),
    ._EVAL_12(widget_1__EVAL_12),
    ._EVAL_13(widget_1__EVAL_13),
    ._EVAL_14(widget_1__EVAL_14),
    ._EVAL_15(widget_1__EVAL_15),
    ._EVAL_16(widget_1__EVAL_16),
    ._EVAL_17(widget_1__EVAL_17),
    ._EVAL_18(widget_1__EVAL_18),
    ._EVAL_19(widget_1__EVAL_19),
    ._EVAL_20(widget_1__EVAL_20),
    ._EVAL_21(widget_1__EVAL_21),
    ._EVAL_22(widget_1__EVAL_22),
    ._EVAL_23(widget_1__EVAL_23),
    ._EVAL_24(widget_1__EVAL_24),
    ._EVAL_25(widget_1__EVAL_25),
    ._EVAL_26(widget_1__EVAL_26),
    ._EVAL_27(widget_1__EVAL_27),
    ._EVAL_28(widget_1__EVAL_28),
    ._EVAL_29(widget_1__EVAL_29),
    ._EVAL_30(widget_1__EVAL_30),
    ._EVAL_31(widget_1__EVAL_31),
    ._EVAL_32(widget_1__EVAL_32)
  );
  SiFive__EVAL_264 filter (
    ._EVAL(filter__EVAL),
    ._EVAL_0(filter__EVAL_0),
    ._EVAL_1(filter__EVAL_1),
    ._EVAL_2(filter__EVAL_2),
    ._EVAL_3(filter__EVAL_3),
    ._EVAL_4(filter__EVAL_4),
    ._EVAL_5(filter__EVAL_5),
    ._EVAL_6(filter__EVAL_6),
    ._EVAL_7(filter__EVAL_7),
    ._EVAL_8(filter__EVAL_8),
    ._EVAL_9(filter__EVAL_9),
    ._EVAL_10(filter__EVAL_10),
    ._EVAL_11(filter__EVAL_11),
    ._EVAL_12(filter__EVAL_12),
    ._EVAL_13(filter__EVAL_13),
    ._EVAL_14(filter__EVAL_14),
    ._EVAL_15(filter__EVAL_15),
    ._EVAL_16(filter__EVAL_16),
    ._EVAL_17(filter__EVAL_17),
    ._EVAL_18(filter__EVAL_18),
    ._EVAL_19(filter__EVAL_19),
    ._EVAL_20(filter__EVAL_20),
    ._EVAL_21(filter__EVAL_21),
    ._EVAL_22(filter__EVAL_22),
    ._EVAL_23(filter__EVAL_23),
    ._EVAL_24(filter__EVAL_24),
    ._EVAL_25(filter__EVAL_25),
    ._EVAL_26(filter__EVAL_26),
    ._EVAL_27(filter__EVAL_27),
    ._EVAL_28(filter__EVAL_28),
    ._EVAL_29(filter__EVAL_29),
    ._EVAL_30(filter__EVAL_30),
    ._EVAL_31(filter__EVAL_31),
    ._EVAL_32(filter__EVAL_32),
    ._EVAL_33(filter__EVAL_33),
    ._EVAL_34(filter__EVAL_34),
    ._EVAL_35(filter__EVAL_35),
    ._EVAL_36(filter__EVAL_36),
    ._EVAL_37(filter__EVAL_37),
    ._EVAL_38(filter__EVAL_38),
    ._EVAL_39(filter__EVAL_39),
    ._EVAL_40(filter__EVAL_40),
    ._EVAL_41(filter__EVAL_41),
    ._EVAL_42(filter__EVAL_42),
    ._EVAL_43(filter__EVAL_43),
    ._EVAL_44(filter__EVAL_44),
    ._EVAL_45(filter__EVAL_45),
    ._EVAL_46(filter__EVAL_46),
    ._EVAL_47(filter__EVAL_47),
    ._EVAL_48(filter__EVAL_48),
    ._EVAL_49(filter__EVAL_49),
    ._EVAL_50(filter__EVAL_50),
    ._EVAL_51(filter__EVAL_51),
    ._EVAL_52(filter__EVAL_52),
    ._EVAL_53(filter__EVAL_53),
    ._EVAL_54(filter__EVAL_54),
    ._EVAL_55(filter__EVAL_55),
    ._EVAL_56(filter__EVAL_56),
    ._EVAL_57(filter__EVAL_57),
    ._EVAL_58(filter__EVAL_58),
    ._EVAL_59(filter__EVAL_59),
    ._EVAL_60(filter__EVAL_60),
    ._EVAL_61(filter__EVAL_61),
    ._EVAL_62(filter__EVAL_62),
    ._EVAL_63(filter__EVAL_63),
    ._EVAL_64(filter__EVAL_64),
    ._EVAL_65(filter__EVAL_65),
    ._EVAL_66(filter__EVAL_66),
    ._EVAL_67(filter__EVAL_67),
    ._EVAL_68(filter__EVAL_68),
    ._EVAL_69(filter__EVAL_69),
    ._EVAL_70(filter__EVAL_70),
    ._EVAL_71(filter__EVAL_71),
    ._EVAL_72(filter__EVAL_72)
  );
  SiFive__EVAL_283 intsink_2 (
    ._EVAL(intsink_2__EVAL),
    ._EVAL_0(intsink_2__EVAL_0),
    ._EVAL_1(intsink_2__EVAL_1)
  );
  SiFive__EVAL_308 FormMicroOps (
    ._EVAL(FormMicroOps__EVAL),
    ._EVAL_0(FormMicroOps__EVAL_0),
    ._EVAL_1(FormMicroOps__EVAL_1),
    ._EVAL_2(FormMicroOps__EVAL_2),
    ._EVAL_3(FormMicroOps__EVAL_3),
    ._EVAL_4(FormMicroOps__EVAL_4),
    ._EVAL_5(FormMicroOps__EVAL_5),
    ._EVAL_6(FormMicroOps__EVAL_6),
    ._EVAL_7(FormMicroOps__EVAL_7),
    ._EVAL_8(FormMicroOps__EVAL_8),
    ._EVAL_9(FormMicroOps__EVAL_9),
    ._EVAL_10(FormMicroOps__EVAL_10),
    ._EVAL_11(FormMicroOps__EVAL_11),
    ._EVAL_12(FormMicroOps__EVAL_12),
    ._EVAL_13(FormMicroOps__EVAL_13),
    ._EVAL_14(FormMicroOps__EVAL_14),
    ._EVAL_15(FormMicroOps__EVAL_15),
    ._EVAL_16(FormMicroOps__EVAL_16),
    ._EVAL_17(FormMicroOps__EVAL_17),
    ._EVAL_18(FormMicroOps__EVAL_18),
    ._EVAL_19(FormMicroOps__EVAL_19),
    ._EVAL_20(FormMicroOps__EVAL_20),
    ._EVAL_21(FormMicroOps__EVAL_21),
    ._EVAL_22(FormMicroOps__EVAL_22),
    ._EVAL_23(FormMicroOps__EVAL_23),
    ._EVAL_24(FormMicroOps__EVAL_24),
    ._EVAL_25(FormMicroOps__EVAL_25),
    ._EVAL_26(FormMicroOps__EVAL_26),
    ._EVAL_27(FormMicroOps__EVAL_27),
    ._EVAL_28(FormMicroOps__EVAL_28),
    ._EVAL_29(FormMicroOps__EVAL_29),
    ._EVAL_30(FormMicroOps__EVAL_30),
    ._EVAL_31(FormMicroOps__EVAL_31),
    ._EVAL_32(FormMicroOps__EVAL_32),
    ._EVAL_33(FormMicroOps__EVAL_33),
    ._EVAL_34(FormMicroOps__EVAL_34),
    ._EVAL_35(FormMicroOps__EVAL_35),
    ._EVAL_36(FormMicroOps__EVAL_36),
    ._EVAL_37(FormMicroOps__EVAL_37),
    ._EVAL_38(FormMicroOps__EVAL_38),
    ._EVAL_39(FormMicroOps__EVAL_39),
    ._EVAL_40(FormMicroOps__EVAL_40),
    ._EVAL_41(FormMicroOps__EVAL_41),
    ._EVAL_42(FormMicroOps__EVAL_42),
    ._EVAL_43(FormMicroOps__EVAL_43),
    ._EVAL_44(FormMicroOps__EVAL_44),
    ._EVAL_45(FormMicroOps__EVAL_45),
    ._EVAL_46(FormMicroOps__EVAL_46),
    ._EVAL_47(FormMicroOps__EVAL_47),
    ._EVAL_48(FormMicroOps__EVAL_48),
    ._EVAL_49(FormMicroOps__EVAL_49),
    ._EVAL_50(FormMicroOps__EVAL_50),
    ._EVAL_51(FormMicroOps__EVAL_51),
    ._EVAL_52(FormMicroOps__EVAL_52),
    ._EVAL_53(FormMicroOps__EVAL_53),
    ._EVAL_54(FormMicroOps__EVAL_54),
    ._EVAL_55(FormMicroOps__EVAL_55),
    ._EVAL_56(FormMicroOps__EVAL_56),
    ._EVAL_57(FormMicroOps__EVAL_57),
    ._EVAL_58(FormMicroOps__EVAL_58),
    ._EVAL_59(FormMicroOps__EVAL_59),
    ._EVAL_60(FormMicroOps__EVAL_60),
    ._EVAL_61(FormMicroOps__EVAL_61),
    ._EVAL_62(FormMicroOps__EVAL_62),
    ._EVAL_63(FormMicroOps__EVAL_63),
    ._EVAL_64(FormMicroOps__EVAL_64),
    ._EVAL_65(FormMicroOps__EVAL_65),
    ._EVAL_66(FormMicroOps__EVAL_66),
    ._EVAL_67(FormMicroOps__EVAL_67),
    ._EVAL_68(FormMicroOps__EVAL_68),
    ._EVAL_69(FormMicroOps__EVAL_69),
    ._EVAL_70(FormMicroOps__EVAL_70),
    ._EVAL_71(FormMicroOps__EVAL_71),
    ._EVAL_72(FormMicroOps__EVAL_72),
    ._EVAL_73(FormMicroOps__EVAL_73),
    ._EVAL_74(FormMicroOps__EVAL_74),
    ._EVAL_75(FormMicroOps__EVAL_75),
    ._EVAL_76(FormMicroOps__EVAL_76),
    ._EVAL_77(FormMicroOps__EVAL_77),
    ._EVAL_78(FormMicroOps__EVAL_78),
    ._EVAL_79(FormMicroOps__EVAL_79),
    ._EVAL_80(FormMicroOps__EVAL_80),
    ._EVAL_81(FormMicroOps__EVAL_81),
    ._EVAL_82(FormMicroOps__EVAL_82),
    ._EVAL_83(FormMicroOps__EVAL_83),
    ._EVAL_84(FormMicroOps__EVAL_84),
    ._EVAL_85(FormMicroOps__EVAL_85),
    ._EVAL_86(FormMicroOps__EVAL_86),
    ._EVAL_87(FormMicroOps__EVAL_87),
    ._EVAL_88(FormMicroOps__EVAL_88),
    ._EVAL_89(FormMicroOps__EVAL_89),
    ._EVAL_90(FormMicroOps__EVAL_90),
    ._EVAL_91(FormMicroOps__EVAL_91),
    ._EVAL_92(FormMicroOps__EVAL_92),
    ._EVAL_93(FormMicroOps__EVAL_93),
    ._EVAL_94(FormMicroOps__EVAL_94),
    ._EVAL_95(FormMicroOps__EVAL_95),
    ._EVAL_96(FormMicroOps__EVAL_96),
    ._EVAL_97(FormMicroOps__EVAL_97),
    ._EVAL_98(FormMicroOps__EVAL_98),
    ._EVAL_99(FormMicroOps__EVAL_99),
    ._EVAL_100(FormMicroOps__EVAL_100),
    ._EVAL_101(FormMicroOps__EVAL_101),
    ._EVAL_102(FormMicroOps__EVAL_102),
    ._EVAL_103(FormMicroOps__EVAL_103),
    ._EVAL_104(FormMicroOps__EVAL_104),
    ._EVAL_105(FormMicroOps__EVAL_105),
    ._EVAL_106(FormMicroOps__EVAL_106),
    ._EVAL_107(FormMicroOps__EVAL_107),
    ._EVAL_108(FormMicroOps__EVAL_108),
    ._EVAL_109(FormMicroOps__EVAL_109),
    ._EVAL_110(FormMicroOps__EVAL_110),
    ._EVAL_111(FormMicroOps__EVAL_111),
    ._EVAL_112(FormMicroOps__EVAL_112),
    ._EVAL_113(FormMicroOps__EVAL_113),
    ._EVAL_114(FormMicroOps__EVAL_114),
    ._EVAL_115(FormMicroOps__EVAL_115),
    ._EVAL_116(FormMicroOps__EVAL_116),
    ._EVAL_117(FormMicroOps__EVAL_117),
    ._EVAL_118(FormMicroOps__EVAL_118),
    ._EVAL_119(FormMicroOps__EVAL_119),
    ._EVAL_120(FormMicroOps__EVAL_120),
    ._EVAL_121(FormMicroOps__EVAL_121),
    ._EVAL_122(FormMicroOps__EVAL_122),
    ._EVAL_123(FormMicroOps__EVAL_123),
    ._EVAL_124(FormMicroOps__EVAL_124),
    ._EVAL_125(FormMicroOps__EVAL_125),
    ._EVAL_126(FormMicroOps__EVAL_126),
    ._EVAL_127(FormMicroOps__EVAL_127),
    ._EVAL_128(FormMicroOps__EVAL_128),
    ._EVAL_129(FormMicroOps__EVAL_129),
    ._EVAL_130(FormMicroOps__EVAL_130),
    ._EVAL_131(FormMicroOps__EVAL_131),
    ._EVAL_132(FormMicroOps__EVAL_132),
    ._EVAL_133(FormMicroOps__EVAL_133),
    ._EVAL_134(FormMicroOps__EVAL_134),
    ._EVAL_135(FormMicroOps__EVAL_135),
    ._EVAL_136(FormMicroOps__EVAL_136),
    ._EVAL_137(FormMicroOps__EVAL_137),
    ._EVAL_138(FormMicroOps__EVAL_138),
    ._EVAL_139(FormMicroOps__EVAL_139),
    ._EVAL_140(FormMicroOps__EVAL_140),
    ._EVAL_141(FormMicroOps__EVAL_141),
    ._EVAL_142(FormMicroOps__EVAL_142),
    ._EVAL_143(FormMicroOps__EVAL_143),
    ._EVAL_144(FormMicroOps__EVAL_144),
    ._EVAL_145(FormMicroOps__EVAL_145),
    ._EVAL_146(FormMicroOps__EVAL_146),
    ._EVAL_147(FormMicroOps__EVAL_147),
    ._EVAL_148(FormMicroOps__EVAL_148),
    ._EVAL_149(FormMicroOps__EVAL_149),
    ._EVAL_150(FormMicroOps__EVAL_150),
    ._EVAL_151(FormMicroOps__EVAL_151),
    ._EVAL_152(FormMicroOps__EVAL_152),
    ._EVAL_153(FormMicroOps__EVAL_153),
    ._EVAL_154(FormMicroOps__EVAL_154),
    ._EVAL_155(FormMicroOps__EVAL_155),
    ._EVAL_156(FormMicroOps__EVAL_156),
    ._EVAL_157(FormMicroOps__EVAL_157),
    ._EVAL_158(FormMicroOps__EVAL_158),
    ._EVAL_159(FormMicroOps__EVAL_159)
  );
  SiFive__EVAL_309 InstructionQueue (
    ._EVAL(InstructionQueue__EVAL),
    ._EVAL_0(InstructionQueue__EVAL_0),
    ._EVAL_1(InstructionQueue__EVAL_1),
    ._EVAL_2(InstructionQueue__EVAL_2),
    ._EVAL_3(InstructionQueue__EVAL_3),
    ._EVAL_4(InstructionQueue__EVAL_4),
    ._EVAL_5(InstructionQueue__EVAL_5),
    ._EVAL_6(InstructionQueue__EVAL_6),
    ._EVAL_7(InstructionQueue__EVAL_7),
    ._EVAL_8(InstructionQueue__EVAL_8),
    ._EVAL_9(InstructionQueue__EVAL_9),
    ._EVAL_10(InstructionQueue__EVAL_10),
    ._EVAL_11(InstructionQueue__EVAL_11),
    ._EVAL_12(InstructionQueue__EVAL_12),
    ._EVAL_13(InstructionQueue__EVAL_13),
    ._EVAL_14(InstructionQueue__EVAL_14),
    ._EVAL_15(InstructionQueue__EVAL_15),
    ._EVAL_16(InstructionQueue__EVAL_16),
    ._EVAL_17(InstructionQueue__EVAL_17),
    ._EVAL_18(InstructionQueue__EVAL_18),
    ._EVAL_19(InstructionQueue__EVAL_19),
    ._EVAL_20(InstructionQueue__EVAL_20),
    ._EVAL_21(InstructionQueue__EVAL_21),
    ._EVAL_22(InstructionQueue__EVAL_22),
    ._EVAL_23(InstructionQueue__EVAL_23),
    ._EVAL_24(InstructionQueue__EVAL_24),
    ._EVAL_25(InstructionQueue__EVAL_25),
    ._EVAL_26(InstructionQueue__EVAL_26),
    ._EVAL_27(InstructionQueue__EVAL_27),
    ._EVAL_28(InstructionQueue__EVAL_28),
    ._EVAL_29(InstructionQueue__EVAL_29),
    ._EVAL_30(InstructionQueue__EVAL_30),
    ._EVAL_31(InstructionQueue__EVAL_31),
    ._EVAL_32(InstructionQueue__EVAL_32),
    ._EVAL_33(InstructionQueue__EVAL_33),
    ._EVAL_34(InstructionQueue__EVAL_34),
    ._EVAL_35(InstructionQueue__EVAL_35),
    ._EVAL_36(InstructionQueue__EVAL_36),
    ._EVAL_37(InstructionQueue__EVAL_37),
    ._EVAL_38(InstructionQueue__EVAL_38),
    ._EVAL_39(InstructionQueue__EVAL_39),
    ._EVAL_40(InstructionQueue__EVAL_40),
    ._EVAL_41(InstructionQueue__EVAL_41),
    ._EVAL_42(InstructionQueue__EVAL_42),
    ._EVAL_43(InstructionQueue__EVAL_43),
    ._EVAL_44(InstructionQueue__EVAL_44),
    ._EVAL_45(InstructionQueue__EVAL_45),
    ._EVAL_46(InstructionQueue__EVAL_46),
    ._EVAL_47(InstructionQueue__EVAL_47),
    ._EVAL_48(InstructionQueue__EVAL_48),
    ._EVAL_49(InstructionQueue__EVAL_49),
    ._EVAL_50(InstructionQueue__EVAL_50),
    ._EVAL_51(InstructionQueue__EVAL_51),
    ._EVAL_52(InstructionQueue__EVAL_52),
    ._EVAL_53(InstructionQueue__EVAL_53),
    ._EVAL_54(InstructionQueue__EVAL_54),
    ._EVAL_55(InstructionQueue__EVAL_55),
    ._EVAL_56(InstructionQueue__EVAL_56),
    ._EVAL_57(InstructionQueue__EVAL_57),
    ._EVAL_58(InstructionQueue__EVAL_58),
    ._EVAL_59(InstructionQueue__EVAL_59),
    ._EVAL_60(InstructionQueue__EVAL_60),
    ._EVAL_61(InstructionQueue__EVAL_61),
    ._EVAL_62(InstructionQueue__EVAL_62),
    ._EVAL_63(InstructionQueue__EVAL_63),
    ._EVAL_64(InstructionQueue__EVAL_64),
    ._EVAL_65(InstructionQueue__EVAL_65),
    ._EVAL_66(InstructionQueue__EVAL_66),
    ._EVAL_67(InstructionQueue__EVAL_67),
    ._EVAL_68(InstructionQueue__EVAL_68),
    ._EVAL_69(InstructionQueue__EVAL_69),
    ._EVAL_70(InstructionQueue__EVAL_70),
    ._EVAL_71(InstructionQueue__EVAL_71),
    ._EVAL_72(InstructionQueue__EVAL_72),
    ._EVAL_73(InstructionQueue__EVAL_73),
    ._EVAL_74(InstructionQueue__EVAL_74),
    ._EVAL_75(InstructionQueue__EVAL_75),
    ._EVAL_76(InstructionQueue__EVAL_76),
    ._EVAL_77(InstructionQueue__EVAL_77),
    ._EVAL_78(InstructionQueue__EVAL_78),
    ._EVAL_79(InstructionQueue__EVAL_79),
    ._EVAL_80(InstructionQueue__EVAL_80),
    ._EVAL_81(InstructionQueue__EVAL_81),
    ._EVAL_82(InstructionQueue__EVAL_82),
    ._EVAL_83(InstructionQueue__EVAL_83),
    ._EVAL_84(InstructionQueue__EVAL_84),
    ._EVAL_85(InstructionQueue__EVAL_85),
    ._EVAL_86(InstructionQueue__EVAL_86),
    ._EVAL_87(InstructionQueue__EVAL_87),
    ._EVAL_88(InstructionQueue__EVAL_88),
    ._EVAL_89(InstructionQueue__EVAL_89),
    ._EVAL_90(InstructionQueue__EVAL_90),
    ._EVAL_91(InstructionQueue__EVAL_91),
    ._EVAL_92(InstructionQueue__EVAL_92),
    ._EVAL_93(InstructionQueue__EVAL_93),
    ._EVAL_94(InstructionQueue__EVAL_94),
    ._EVAL_95(InstructionQueue__EVAL_95),
    ._EVAL_96(InstructionQueue__EVAL_96),
    ._EVAL_97(InstructionQueue__EVAL_97),
    ._EVAL_98(InstructionQueue__EVAL_98),
    ._EVAL_99(InstructionQueue__EVAL_99),
    ._EVAL_100(InstructionQueue__EVAL_100),
    ._EVAL_101(InstructionQueue__EVAL_101),
    ._EVAL_102(InstructionQueue__EVAL_102),
    ._EVAL_103(InstructionQueue__EVAL_103),
    ._EVAL_104(InstructionQueue__EVAL_104),
    ._EVAL_105(InstructionQueue__EVAL_105),
    ._EVAL_106(InstructionQueue__EVAL_106),
    ._EVAL_107(InstructionQueue__EVAL_107),
    ._EVAL_108(InstructionQueue__EVAL_108),
    ._EVAL_109(InstructionQueue__EVAL_109),
    ._EVAL_110(InstructionQueue__EVAL_110),
    ._EVAL_111(InstructionQueue__EVAL_111),
    ._EVAL_112(InstructionQueue__EVAL_112),
    ._EVAL_113(InstructionQueue__EVAL_113),
    ._EVAL_114(InstructionQueue__EVAL_114),
    ._EVAL_115(InstructionQueue__EVAL_115),
    ._EVAL_116(InstructionQueue__EVAL_116),
    ._EVAL_117(InstructionQueue__EVAL_117),
    ._EVAL_118(InstructionQueue__EVAL_118),
    ._EVAL_119(InstructionQueue__EVAL_119),
    ._EVAL_120(InstructionQueue__EVAL_120),
    ._EVAL_121(InstructionQueue__EVAL_121),
    ._EVAL_122(InstructionQueue__EVAL_122),
    ._EVAL_123(InstructionQueue__EVAL_123),
    ._EVAL_124(InstructionQueue__EVAL_124),
    ._EVAL_125(InstructionQueue__EVAL_125),
    ._EVAL_126(InstructionQueue__EVAL_126),
    ._EVAL_127(InstructionQueue__EVAL_127),
    ._EVAL_128(InstructionQueue__EVAL_128),
    ._EVAL_129(InstructionQueue__EVAL_129),
    ._EVAL_130(InstructionQueue__EVAL_130),
    ._EVAL_131(InstructionQueue__EVAL_131),
    ._EVAL_132(InstructionQueue__EVAL_132),
    ._EVAL_133(InstructionQueue__EVAL_133),
    ._EVAL_134(InstructionQueue__EVAL_134),
    ._EVAL_135(InstructionQueue__EVAL_135),
    ._EVAL_136(InstructionQueue__EVAL_136),
    ._EVAL_137(InstructionQueue__EVAL_137),
    ._EVAL_138(InstructionQueue__EVAL_138),
    ._EVAL_139(InstructionQueue__EVAL_139),
    ._EVAL_140(InstructionQueue__EVAL_140),
    ._EVAL_141(InstructionQueue__EVAL_141),
    ._EVAL_142(InstructionQueue__EVAL_142),
    ._EVAL_143(InstructionQueue__EVAL_143),
    ._EVAL_144(InstructionQueue__EVAL_144),
    ._EVAL_145(InstructionQueue__EVAL_145),
    ._EVAL_146(InstructionQueue__EVAL_146),
    ._EVAL_147(InstructionQueue__EVAL_147),
    ._EVAL_148(InstructionQueue__EVAL_148),
    ._EVAL_149(InstructionQueue__EVAL_149),
    ._EVAL_150(InstructionQueue__EVAL_150),
    ._EVAL_151(InstructionQueue__EVAL_151),
    ._EVAL_152(InstructionQueue__EVAL_152),
    ._EVAL_153(InstructionQueue__EVAL_153),
    ._EVAL_154(InstructionQueue__EVAL_154),
    ._EVAL_155(InstructionQueue__EVAL_155),
    ._EVAL_156(InstructionQueue__EVAL_156),
    ._EVAL_157(InstructionQueue__EVAL_157),
    ._EVAL_158(InstructionQueue__EVAL_158),
    ._EVAL_159(InstructionQueue__EVAL_159),
    ._EVAL_160(InstructionQueue__EVAL_160),
    ._EVAL_161(InstructionQueue__EVAL_161),
    ._EVAL_162(InstructionQueue__EVAL_162),
    ._EVAL_163(InstructionQueue__EVAL_163),
    ._EVAL_164(InstructionQueue__EVAL_164),
    ._EVAL_165(InstructionQueue__EVAL_165),
    ._EVAL_166(InstructionQueue__EVAL_166),
    ._EVAL_167(InstructionQueue__EVAL_167),
    ._EVAL_168(InstructionQueue__EVAL_168),
    ._EVAL_169(InstructionQueue__EVAL_169),
    ._EVAL_170(InstructionQueue__EVAL_170),
    ._EVAL_171(InstructionQueue__EVAL_171),
    ._EVAL_172(InstructionQueue__EVAL_172),
    ._EVAL_173(InstructionQueue__EVAL_173),
    ._EVAL_174(InstructionQueue__EVAL_174),
    ._EVAL_175(InstructionQueue__EVAL_175),
    ._EVAL_176(InstructionQueue__EVAL_176),
    ._EVAL_177(InstructionQueue__EVAL_177),
    ._EVAL_178(InstructionQueue__EVAL_178),
    ._EVAL_179(InstructionQueue__EVAL_179),
    ._EVAL_180(InstructionQueue__EVAL_180),
    ._EVAL_181(InstructionQueue__EVAL_181),
    ._EVAL_182(InstructionQueue__EVAL_182),
    ._EVAL_183(InstructionQueue__EVAL_183),
    ._EVAL_184(InstructionQueue__EVAL_184),
    ._EVAL_185(InstructionQueue__EVAL_185)
  );
  SiFive__EVAL_226 tlSlaveXbar (
    ._EVAL(tlSlaveXbar__EVAL),
    ._EVAL_0(tlSlaveXbar__EVAL_0),
    ._EVAL_1(tlSlaveXbar__EVAL_1),
    ._EVAL_2(tlSlaveXbar__EVAL_2),
    ._EVAL_3(tlSlaveXbar__EVAL_3),
    ._EVAL_4(tlSlaveXbar__EVAL_4),
    ._EVAL_5(tlSlaveXbar__EVAL_5),
    ._EVAL_6(tlSlaveXbar__EVAL_6),
    ._EVAL_7(tlSlaveXbar__EVAL_7),
    ._EVAL_8(tlSlaveXbar__EVAL_8),
    ._EVAL_9(tlSlaveXbar__EVAL_9),
    ._EVAL_10(tlSlaveXbar__EVAL_10),
    ._EVAL_11(tlSlaveXbar__EVAL_11),
    ._EVAL_12(tlSlaveXbar__EVAL_12),
    ._EVAL_13(tlSlaveXbar__EVAL_13),
    ._EVAL_14(tlSlaveXbar__EVAL_14),
    ._EVAL_15(tlSlaveXbar__EVAL_15),
    ._EVAL_16(tlSlaveXbar__EVAL_16),
    ._EVAL_17(tlSlaveXbar__EVAL_17),
    ._EVAL_18(tlSlaveXbar__EVAL_18),
    ._EVAL_19(tlSlaveXbar__EVAL_19),
    ._EVAL_20(tlSlaveXbar__EVAL_20),
    ._EVAL_21(tlSlaveXbar__EVAL_21),
    ._EVAL_22(tlSlaveXbar__EVAL_22),
    ._EVAL_23(tlSlaveXbar__EVAL_23),
    ._EVAL_24(tlSlaveXbar__EVAL_24),
    ._EVAL_25(tlSlaveXbar__EVAL_25),
    ._EVAL_26(tlSlaveXbar__EVAL_26),
    ._EVAL_27(tlSlaveXbar__EVAL_27),
    ._EVAL_28(tlSlaveXbar__EVAL_28),
    ._EVAL_29(tlSlaveXbar__EVAL_29),
    ._EVAL_30(tlSlaveXbar__EVAL_30),
    ._EVAL_31(tlSlaveXbar__EVAL_31),
    ._EVAL_32(tlSlaveXbar__EVAL_32),
    ._EVAL_33(tlSlaveXbar__EVAL_33),
    ._EVAL_34(tlSlaveXbar__EVAL_34),
    ._EVAL_35(tlSlaveXbar__EVAL_35),
    ._EVAL_36(tlSlaveXbar__EVAL_36),
    ._EVAL_37(tlSlaveXbar__EVAL_37),
    ._EVAL_38(tlSlaveXbar__EVAL_38),
    ._EVAL_39(tlSlaveXbar__EVAL_39),
    ._EVAL_40(tlSlaveXbar__EVAL_40),
    ._EVAL_41(tlSlaveXbar__EVAL_41),
    ._EVAL_42(tlSlaveXbar__EVAL_42),
    ._EVAL_43(tlSlaveXbar__EVAL_43),
    ._EVAL_44(tlSlaveXbar__EVAL_44),
    ._EVAL_45(tlSlaveXbar__EVAL_45),
    ._EVAL_46(tlSlaveXbar__EVAL_46),
    ._EVAL_47(tlSlaveXbar__EVAL_47),
    ._EVAL_48(tlSlaveXbar__EVAL_48),
    ._EVAL_49(tlSlaveXbar__EVAL_49),
    ._EVAL_50(tlSlaveXbar__EVAL_50)
  );
  SiFive__EVAL_266 buffer_2 (
    ._EVAL(buffer_2__EVAL),
    ._EVAL_0(buffer_2__EVAL_0),
    ._EVAL_1(buffer_2__EVAL_1),
    ._EVAL_2(buffer_2__EVAL_2),
    ._EVAL_3(buffer_2__EVAL_3),
    ._EVAL_4(buffer_2__EVAL_4),
    ._EVAL_5(buffer_2__EVAL_5),
    ._EVAL_6(buffer_2__EVAL_6),
    ._EVAL_7(buffer_2__EVAL_7),
    ._EVAL_8(buffer_2__EVAL_8),
    ._EVAL_9(buffer_2__EVAL_9),
    ._EVAL_10(buffer_2__EVAL_10),
    ._EVAL_11(buffer_2__EVAL_11),
    ._EVAL_12(buffer_2__EVAL_12),
    ._EVAL_13(buffer_2__EVAL_13),
    ._EVAL_14(buffer_2__EVAL_14),
    ._EVAL_15(buffer_2__EVAL_15),
    ._EVAL_16(buffer_2__EVAL_16),
    ._EVAL_17(buffer_2__EVAL_17),
    ._EVAL_18(buffer_2__EVAL_18),
    ._EVAL_19(buffer_2__EVAL_19),
    ._EVAL_20(buffer_2__EVAL_20),
    ._EVAL_21(buffer_2__EVAL_21),
    ._EVAL_22(buffer_2__EVAL_22),
    ._EVAL_23(buffer_2__EVAL_23),
    ._EVAL_24(buffer_2__EVAL_24),
    ._EVAL_25(buffer_2__EVAL_25),
    ._EVAL_26(buffer_2__EVAL_26),
    ._EVAL_27(buffer_2__EVAL_27),
    ._EVAL_28(buffer_2__EVAL_28),
    ._EVAL_29(buffer_2__EVAL_29),
    ._EVAL_30(buffer_2__EVAL_30),
    ._EVAL_31(buffer_2__EVAL_31),
    ._EVAL_32(buffer_2__EVAL_32),
    ._EVAL_33(buffer_2__EVAL_33),
    ._EVAL_34(buffer_2__EVAL_34),
    ._EVAL_35(buffer_2__EVAL_35),
    ._EVAL_36(buffer_2__EVAL_36),
    ._EVAL_37(buffer_2__EVAL_37),
    ._EVAL_38(buffer_2__EVAL_38),
    ._EVAL_39(buffer_2__EVAL_39),
    ._EVAL_40(buffer_2__EVAL_40),
    ._EVAL_41(buffer_2__EVAL_41),
    ._EVAL_42(buffer_2__EVAL_42),
    ._EVAL_43(buffer_2__EVAL_43),
    ._EVAL_44(buffer_2__EVAL_44),
    ._EVAL_45(buffer_2__EVAL_45),
    ._EVAL_46(buffer_2__EVAL_46),
    ._EVAL_47(buffer_2__EVAL_47),
    ._EVAL_48(buffer_2__EVAL_48),
    ._EVAL_49(buffer_2__EVAL_49),
    ._EVAL_50(buffer_2__EVAL_50),
    ._EVAL_51(buffer_2__EVAL_51),
    ._EVAL_52(buffer_2__EVAL_52),
    ._EVAL_53(buffer_2__EVAL_53),
    ._EVAL_54(buffer_2__EVAL_54),
    ._EVAL_55(buffer_2__EVAL_55),
    ._EVAL_56(buffer_2__EVAL_56),
    ._EVAL_57(buffer_2__EVAL_57),
    ._EVAL_58(buffer_2__EVAL_58),
    ._EVAL_59(buffer_2__EVAL_59),
    ._EVAL_60(buffer_2__EVAL_60),
    ._EVAL_61(buffer_2__EVAL_61),
    ._EVAL_62(buffer_2__EVAL_62),
    ._EVAL_63(buffer_2__EVAL_63),
    ._EVAL_64(buffer_2__EVAL_64),
    ._EVAL_65(buffer_2__EVAL_65),
    ._EVAL_66(buffer_2__EVAL_66),
    ._EVAL_67(buffer_2__EVAL_67),
    ._EVAL_68(buffer_2__EVAL_68),
    ._EVAL_69(buffer_2__EVAL_69),
    ._EVAL_70(buffer_2__EVAL_70),
    ._EVAL_71(buffer_2__EVAL_71),
    ._EVAL_72(buffer_2__EVAL_72)
  );
  SiFive__EVAL_251 buffer_1 (
    ._EVAL(buffer_1__EVAL),
    ._EVAL_0(buffer_1__EVAL_0),
    ._EVAL_1(buffer_1__EVAL_1),
    ._EVAL_2(buffer_1__EVAL_2),
    ._EVAL_3(buffer_1__EVAL_3),
    ._EVAL_4(buffer_1__EVAL_4),
    ._EVAL_5(buffer_1__EVAL_5),
    ._EVAL_6(buffer_1__EVAL_6),
    ._EVAL_7(buffer_1__EVAL_7),
    ._EVAL_8(buffer_1__EVAL_8),
    ._EVAL_9(buffer_1__EVAL_9),
    ._EVAL_10(buffer_1__EVAL_10),
    ._EVAL_11(buffer_1__EVAL_11),
    ._EVAL_12(buffer_1__EVAL_12),
    ._EVAL_13(buffer_1__EVAL_13),
    ._EVAL_14(buffer_1__EVAL_14),
    ._EVAL_15(buffer_1__EVAL_15),
    ._EVAL_16(buffer_1__EVAL_16),
    ._EVAL_17(buffer_1__EVAL_17),
    ._EVAL_18(buffer_1__EVAL_18),
    ._EVAL_19(buffer_1__EVAL_19),
    ._EVAL_20(buffer_1__EVAL_20),
    ._EVAL_21(buffer_1__EVAL_21),
    ._EVAL_22(buffer_1__EVAL_22),
    ._EVAL_23(buffer_1__EVAL_23),
    ._EVAL_24(buffer_1__EVAL_24),
    ._EVAL_25(buffer_1__EVAL_25),
    ._EVAL_26(buffer_1__EVAL_26),
    ._EVAL_27(buffer_1__EVAL_27),
    ._EVAL_28(buffer_1__EVAL_28),
    ._EVAL_29(buffer_1__EVAL_29),
    ._EVAL_30(buffer_1__EVAL_30),
    ._EVAL_31(buffer_1__EVAL_31),
    ._EVAL_32(buffer_1__EVAL_32)
  );
  SiFive__EVAL_284 dcacheArb (
    ._EVAL(dcacheArb__EVAL),
    ._EVAL_0(dcacheArb__EVAL_0),
    ._EVAL_1(dcacheArb__EVAL_1),
    ._EVAL_2(dcacheArb__EVAL_2),
    ._EVAL_3(dcacheArb__EVAL_3),
    ._EVAL_4(dcacheArb__EVAL_4),
    ._EVAL_5(dcacheArb__EVAL_5),
    ._EVAL_6(dcacheArb__EVAL_6),
    ._EVAL_7(dcacheArb__EVAL_7),
    ._EVAL_8(dcacheArb__EVAL_8),
    ._EVAL_9(dcacheArb__EVAL_9),
    ._EVAL_10(dcacheArb__EVAL_10),
    ._EVAL_11(dcacheArb__EVAL_11),
    ._EVAL_12(dcacheArb__EVAL_12),
    ._EVAL_13(dcacheArb__EVAL_13),
    ._EVAL_14(dcacheArb__EVAL_14),
    ._EVAL_15(dcacheArb__EVAL_15),
    ._EVAL_16(dcacheArb__EVAL_16),
    ._EVAL_17(dcacheArb__EVAL_17),
    ._EVAL_18(dcacheArb__EVAL_18),
    ._EVAL_19(dcacheArb__EVAL_19),
    ._EVAL_20(dcacheArb__EVAL_20),
    ._EVAL_21(dcacheArb__EVAL_21),
    ._EVAL_22(dcacheArb__EVAL_22),
    ._EVAL_23(dcacheArb__EVAL_23),
    ._EVAL_24(dcacheArb__EVAL_24),
    ._EVAL_25(dcacheArb__EVAL_25),
    ._EVAL_26(dcacheArb__EVAL_26),
    ._EVAL_27(dcacheArb__EVAL_27),
    ._EVAL_28(dcacheArb__EVAL_28),
    ._EVAL_29(dcacheArb__EVAL_29),
    ._EVAL_30(dcacheArb__EVAL_30),
    ._EVAL_31(dcacheArb__EVAL_31),
    ._EVAL_32(dcacheArb__EVAL_32),
    ._EVAL_33(dcacheArb__EVAL_33),
    ._EVAL_34(dcacheArb__EVAL_34),
    ._EVAL_35(dcacheArb__EVAL_35),
    ._EVAL_36(dcacheArb__EVAL_36),
    ._EVAL_37(dcacheArb__EVAL_37),
    ._EVAL_38(dcacheArb__EVAL_38),
    ._EVAL_39(dcacheArb__EVAL_39),
    ._EVAL_40(dcacheArb__EVAL_40),
    ._EVAL_41(dcacheArb__EVAL_41),
    ._EVAL_42(dcacheArb__EVAL_42),
    ._EVAL_43(dcacheArb__EVAL_43),
    ._EVAL_44(dcacheArb__EVAL_44),
    ._EVAL_45(dcacheArb__EVAL_45),
    ._EVAL_46(dcacheArb__EVAL_46),
    ._EVAL_47(dcacheArb__EVAL_47),
    ._EVAL_48(dcacheArb__EVAL_48),
    ._EVAL_49(dcacheArb__EVAL_49),
    ._EVAL_50(dcacheArb__EVAL_50),
    ._EVAL_51(dcacheArb__EVAL_51),
    ._EVAL_52(dcacheArb__EVAL_52),
    ._EVAL_53(dcacheArb__EVAL_53),
    ._EVAL_54(dcacheArb__EVAL_54),
    ._EVAL_55(dcacheArb__EVAL_55),
    ._EVAL_56(dcacheArb__EVAL_56),
    ._EVAL_57(dcacheArb__EVAL_57),
    ._EVAL_58(dcacheArb__EVAL_58),
    ._EVAL_59(dcacheArb__EVAL_59),
    ._EVAL_60(dcacheArb__EVAL_60),
    ._EVAL_61(dcacheArb__EVAL_61),
    ._EVAL_62(dcacheArb__EVAL_62),
    ._EVAL_63(dcacheArb__EVAL_63),
    ._EVAL_64(dcacheArb__EVAL_64),
    ._EVAL_65(dcacheArb__EVAL_65),
    ._EVAL_66(dcacheArb__EVAL_66),
    ._EVAL_67(dcacheArb__EVAL_67),
    ._EVAL_68(dcacheArb__EVAL_68),
    ._EVAL_69(dcacheArb__EVAL_69),
    ._EVAL_70(dcacheArb__EVAL_70),
    ._EVAL_71(dcacheArb__EVAL_71),
    ._EVAL_72(dcacheArb__EVAL_72),
    ._EVAL_73(dcacheArb__EVAL_73),
    ._EVAL_74(dcacheArb__EVAL_74),
    ._EVAL_75(dcacheArb__EVAL_75),
    ._EVAL_76(dcacheArb__EVAL_76),
    ._EVAL_77(dcacheArb__EVAL_77),
    ._EVAL_78(dcacheArb__EVAL_78),
    ._EVAL_79(dcacheArb__EVAL_79),
    ._EVAL_80(dcacheArb__EVAL_80),
    ._EVAL_81(dcacheArb__EVAL_81),
    ._EVAL_82(dcacheArb__EVAL_82),
    ._EVAL_83(dcacheArb__EVAL_83),
    ._EVAL_84(dcacheArb__EVAL_84),
    ._EVAL_85(dcacheArb__EVAL_85),
    ._EVAL_86(dcacheArb__EVAL_86),
    ._EVAL_87(dcacheArb__EVAL_87),
    ._EVAL_88(dcacheArb__EVAL_88),
    ._EVAL_89(dcacheArb__EVAL_89),
    ._EVAL_90(dcacheArb__EVAL_90)
  );
  SiFive__EVAL_274 buffer_3 (
    ._EVAL(buffer_3__EVAL),
    ._EVAL_0(buffer_3__EVAL_0),
    ._EVAL_1(buffer_3__EVAL_1),
    ._EVAL_2(buffer_3__EVAL_2),
    ._EVAL_3(buffer_3__EVAL_3),
    ._EVAL_4(buffer_3__EVAL_4),
    ._EVAL_5(buffer_3__EVAL_5),
    ._EVAL_6(buffer_3__EVAL_6),
    ._EVAL_7(buffer_3__EVAL_7),
    ._EVAL_8(buffer_3__EVAL_8),
    ._EVAL_9(buffer_3__EVAL_9),
    ._EVAL_10(buffer_3__EVAL_10),
    ._EVAL_11(buffer_3__EVAL_11),
    ._EVAL_12(buffer_3__EVAL_12),
    ._EVAL_13(buffer_3__EVAL_13),
    ._EVAL_14(buffer_3__EVAL_14),
    ._EVAL_15(buffer_3__EVAL_15),
    ._EVAL_16(buffer_3__EVAL_16),
    ._EVAL_17(buffer_3__EVAL_17),
    ._EVAL_18(buffer_3__EVAL_18),
    ._EVAL_19(buffer_3__EVAL_19),
    ._EVAL_20(buffer_3__EVAL_20),
    ._EVAL_21(buffer_3__EVAL_21),
    ._EVAL_22(buffer_3__EVAL_22),
    ._EVAL_23(buffer_3__EVAL_23),
    ._EVAL_24(buffer_3__EVAL_24),
    ._EVAL_25(buffer_3__EVAL_25),
    ._EVAL_26(buffer_3__EVAL_26),
    ._EVAL_27(buffer_3__EVAL_27),
    ._EVAL_28(buffer_3__EVAL_28),
    ._EVAL_29(buffer_3__EVAL_29),
    ._EVAL_30(buffer_3__EVAL_30),
    ._EVAL_31(buffer_3__EVAL_31),
    ._EVAL_32(buffer_3__EVAL_32),
    ._EVAL_33(buffer_3__EVAL_33),
    ._EVAL_34(buffer_3__EVAL_34),
    ._EVAL_35(buffer_3__EVAL_35),
    ._EVAL_36(buffer_3__EVAL_36),
    ._EVAL_37(buffer_3__EVAL_37),
    ._EVAL_38(buffer_3__EVAL_38)
  );
  SiFive__EVAL_253 coreXbar (
    ._EVAL(coreXbar__EVAL),
    ._EVAL_0(coreXbar__EVAL_0),
    ._EVAL_1(coreXbar__EVAL_1),
    ._EVAL_2(coreXbar__EVAL_2),
    ._EVAL_3(coreXbar__EVAL_3),
    ._EVAL_4(coreXbar__EVAL_4),
    ._EVAL_5(coreXbar__EVAL_5),
    ._EVAL_6(coreXbar__EVAL_6),
    ._EVAL_7(coreXbar__EVAL_7),
    ._EVAL_8(coreXbar__EVAL_8),
    ._EVAL_9(coreXbar__EVAL_9),
    ._EVAL_10(coreXbar__EVAL_10),
    ._EVAL_11(coreXbar__EVAL_11),
    ._EVAL_12(coreXbar__EVAL_12),
    ._EVAL_13(coreXbar__EVAL_13),
    ._EVAL_14(coreXbar__EVAL_14),
    ._EVAL_15(coreXbar__EVAL_15),
    ._EVAL_16(coreXbar__EVAL_16),
    ._EVAL_17(coreXbar__EVAL_17),
    ._EVAL_18(coreXbar__EVAL_18),
    ._EVAL_19(coreXbar__EVAL_19),
    ._EVAL_20(coreXbar__EVAL_20),
    ._EVAL_21(coreXbar__EVAL_21),
    ._EVAL_22(coreXbar__EVAL_22),
    ._EVAL_23(coreXbar__EVAL_23),
    ._EVAL_24(coreXbar__EVAL_24),
    ._EVAL_25(coreXbar__EVAL_25),
    ._EVAL_26(coreXbar__EVAL_26),
    ._EVAL_27(coreXbar__EVAL_27),
    ._EVAL_28(coreXbar__EVAL_28),
    ._EVAL_29(coreXbar__EVAL_29),
    ._EVAL_30(coreXbar__EVAL_30),
    ._EVAL_31(coreXbar__EVAL_31),
    ._EVAL_32(coreXbar__EVAL_32),
    ._EVAL_33(coreXbar__EVAL_33),
    ._EVAL_34(coreXbar__EVAL_34),
    ._EVAL_35(coreXbar__EVAL_35),
    ._EVAL_36(coreXbar__EVAL_36),
    ._EVAL_37(coreXbar__EVAL_37),
    ._EVAL_38(coreXbar__EVAL_38),
    ._EVAL_39(coreXbar__EVAL_39),
    ._EVAL_40(coreXbar__EVAL_40),
    ._EVAL_41(coreXbar__EVAL_41),
    ._EVAL_42(coreXbar__EVAL_42),
    ._EVAL_43(coreXbar__EVAL_43),
    ._EVAL_44(coreXbar__EVAL_44),
    ._EVAL_45(coreXbar__EVAL_45),
    ._EVAL_46(coreXbar__EVAL_46),
    ._EVAL_47(coreXbar__EVAL_47),
    ._EVAL_48(coreXbar__EVAL_48),
    ._EVAL_49(coreXbar__EVAL_49),
    ._EVAL_50(coreXbar__EVAL_50),
    ._EVAL_51(coreXbar__EVAL_51),
    ._EVAL_52(coreXbar__EVAL_52),
    ._EVAL_53(coreXbar__EVAL_53),
    ._EVAL_54(coreXbar__EVAL_54),
    ._EVAL_55(coreXbar__EVAL_55),
    ._EVAL_56(coreXbar__EVAL_56),
    ._EVAL_57(coreXbar__EVAL_57),
    ._EVAL_58(coreXbar__EVAL_58),
    ._EVAL_59(coreXbar__EVAL_59),
    ._EVAL_60(coreXbar__EVAL_60),
    ._EVAL_61(coreXbar__EVAL_61),
    ._EVAL_62(coreXbar__EVAL_62),
    ._EVAL_63(coreXbar__EVAL_63),
    ._EVAL_64(coreXbar__EVAL_64),
    ._EVAL_65(coreXbar__EVAL_65),
    ._EVAL_66(coreXbar__EVAL_66),
    ._EVAL_67(coreXbar__EVAL_67),
    ._EVAL_68(coreXbar__EVAL_68),
    ._EVAL_69(coreXbar__EVAL_69),
    ._EVAL_70(coreXbar__EVAL_70),
    ._EVAL_71(coreXbar__EVAL_71),
    ._EVAL_72(coreXbar__EVAL_72),
    ._EVAL_73(coreXbar__EVAL_73),
    ._EVAL_74(coreXbar__EVAL_74),
    ._EVAL_75(coreXbar__EVAL_75),
    ._EVAL_76(coreXbar__EVAL_76),
    ._EVAL_77(coreXbar__EVAL_77),
    ._EVAL_78(coreXbar__EVAL_78),
    ._EVAL_79(coreXbar__EVAL_79),
    ._EVAL_80(coreXbar__EVAL_80),
    ._EVAL_81(coreXbar__EVAL_81),
    ._EVAL_82(coreXbar__EVAL_82),
    ._EVAL_83(coreXbar__EVAL_83),
    ._EVAL_84(coreXbar__EVAL_84),
    ._EVAL_85(coreXbar__EVAL_85),
    ._EVAL_86(coreXbar__EVAL_86),
    ._EVAL_87(coreXbar__EVAL_87),
    ._EVAL_88(coreXbar__EVAL_88)
  );
  SiFive__EVAL_227 intXbar (
    ._EVAL(intXbar__EVAL),
    ._EVAL_0(intXbar__EVAL_0),
    ._EVAL_1(intXbar__EVAL_1),
    ._EVAL_2(intXbar__EVAL_2),
    ._EVAL_3(intXbar__EVAL_3),
    ._EVAL_4(intXbar__EVAL_4),
    ._EVAL_5(intXbar__EVAL_5),
    ._EVAL_6(intXbar__EVAL_6)
  );
  SiFive__EVAL_225 tlMasterXbar (
    ._EVAL(tlMasterXbar__EVAL),
    ._EVAL_0(tlMasterXbar__EVAL_0),
    ._EVAL_1(tlMasterXbar__EVAL_1),
    ._EVAL_2(tlMasterXbar__EVAL_2),
    ._EVAL_3(tlMasterXbar__EVAL_3),
    ._EVAL_4(tlMasterXbar__EVAL_4),
    ._EVAL_5(tlMasterXbar__EVAL_5),
    ._EVAL_6(tlMasterXbar__EVAL_6),
    ._EVAL_7(tlMasterXbar__EVAL_7),
    ._EVAL_8(tlMasterXbar__EVAL_8),
    ._EVAL_9(tlMasterXbar__EVAL_9),
    ._EVAL_10(tlMasterXbar__EVAL_10),
    ._EVAL_11(tlMasterXbar__EVAL_11),
    ._EVAL_12(tlMasterXbar__EVAL_12),
    ._EVAL_13(tlMasterXbar__EVAL_13),
    ._EVAL_14(tlMasterXbar__EVAL_14),
    ._EVAL_15(tlMasterXbar__EVAL_15),
    ._EVAL_16(tlMasterXbar__EVAL_16),
    ._EVAL_17(tlMasterXbar__EVAL_17),
    ._EVAL_18(tlMasterXbar__EVAL_18),
    ._EVAL_19(tlMasterXbar__EVAL_19),
    ._EVAL_20(tlMasterXbar__EVAL_20),
    ._EVAL_21(tlMasterXbar__EVAL_21),
    ._EVAL_22(tlMasterXbar__EVAL_22),
    ._EVAL_23(tlMasterXbar__EVAL_23),
    ._EVAL_24(tlMasterXbar__EVAL_24),
    ._EVAL_25(tlMasterXbar__EVAL_25),
    ._EVAL_26(tlMasterXbar__EVAL_26),
    ._EVAL_27(tlMasterXbar__EVAL_27),
    ._EVAL_28(tlMasterXbar__EVAL_28),
    ._EVAL_29(tlMasterXbar__EVAL_29),
    ._EVAL_30(tlMasterXbar__EVAL_30),
    ._EVAL_31(tlMasterXbar__EVAL_31),
    ._EVAL_32(tlMasterXbar__EVAL_32),
    ._EVAL_33(tlMasterXbar__EVAL_33),
    ._EVAL_34(tlMasterXbar__EVAL_34),
    ._EVAL_35(tlMasterXbar__EVAL_35),
    ._EVAL_36(tlMasterXbar__EVAL_36),
    ._EVAL_37(tlMasterXbar__EVAL_37),
    ._EVAL_38(tlMasterXbar__EVAL_38),
    ._EVAL_39(tlMasterXbar__EVAL_39),
    ._EVAL_40(tlMasterXbar__EVAL_40),
    ._EVAL_41(tlMasterXbar__EVAL_41),
    ._EVAL_42(tlMasterXbar__EVAL_42),
    ._EVAL_43(tlMasterXbar__EVAL_43),
    ._EVAL_44(tlMasterXbar__EVAL_44),
    ._EVAL_45(tlMasterXbar__EVAL_45),
    ._EVAL_46(tlMasterXbar__EVAL_46),
    ._EVAL_47(tlMasterXbar__EVAL_47),
    ._EVAL_48(tlMasterXbar__EVAL_48),
    ._EVAL_49(tlMasterXbar__EVAL_49),
    ._EVAL_50(tlMasterXbar__EVAL_50),
    ._EVAL_51(tlMasterXbar__EVAL_51),
    ._EVAL_52(tlMasterXbar__EVAL_52),
    ._EVAL_53(tlMasterXbar__EVAL_53),
    ._EVAL_54(tlMasterXbar__EVAL_54),
    ._EVAL_55(tlMasterXbar__EVAL_55),
    ._EVAL_56(tlMasterXbar__EVAL_56),
    ._EVAL_57(tlMasterXbar__EVAL_57),
    ._EVAL_58(tlMasterXbar__EVAL_58),
    ._EVAL_59(tlMasterXbar__EVAL_59),
    ._EVAL_60(tlMasterXbar__EVAL_60),
    ._EVAL_61(tlMasterXbar__EVAL_61),
    ._EVAL_62(tlMasterXbar__EVAL_62),
    ._EVAL_63(tlMasterXbar__EVAL_63),
    ._EVAL_64(tlMasterXbar__EVAL_64),
    ._EVAL_65(tlMasterXbar__EVAL_65),
    ._EVAL_66(tlMasterXbar__EVAL_66),
    ._EVAL_67(tlMasterXbar__EVAL_67),
    ._EVAL_68(tlMasterXbar__EVAL_68),
    ._EVAL_69(tlMasterXbar__EVAL_69),
    ._EVAL_70(tlMasterXbar__EVAL_70),
    ._EVAL_71(tlMasterXbar__EVAL_71),
    ._EVAL_72(tlMasterXbar__EVAL_72),
    ._EVAL_73(tlMasterXbar__EVAL_73),
    ._EVAL_74(tlMasterXbar__EVAL_74),
    ._EVAL_75(tlMasterXbar__EVAL_75),
    ._EVAL_76(tlMasterXbar__EVAL_76),
    ._EVAL_77(tlMasterXbar__EVAL_77),
    ._EVAL_78(tlMasterXbar__EVAL_78),
    ._EVAL_79(tlMasterXbar__EVAL_79),
    ._EVAL_80(tlMasterXbar__EVAL_80),
    ._EVAL_81(tlMasterXbar__EVAL_81),
    ._EVAL_82(tlMasterXbar__EVAL_82),
    ._EVAL_83(tlMasterXbar__EVAL_83)
  );
  SiFive__EVAL_273 rsource (
    ._EVAL(rsource__EVAL),
    ._EVAL_0(rsource__EVAL_0),
    ._EVAL_1(rsource__EVAL_1),
    ._EVAL_2(rsource__EVAL_2),
    ._EVAL_3(rsource__EVAL_3),
    ._EVAL_4(rsource__EVAL_4),
    ._EVAL_5(rsource__EVAL_5),
    ._EVAL_6(rsource__EVAL_6),
    ._EVAL_7(rsource__EVAL_7),
    ._EVAL_8(rsource__EVAL_8),
    ._EVAL_9(rsource__EVAL_9),
    ._EVAL_10(rsource__EVAL_10),
    ._EVAL_11(rsource__EVAL_11),
    ._EVAL_12(rsource__EVAL_12),
    ._EVAL_13(rsource__EVAL_13),
    ._EVAL_14(rsource__EVAL_14),
    ._EVAL_15(rsource__EVAL_15),
    ._EVAL_16(rsource__EVAL_16),
    ._EVAL_17(rsource__EVAL_17),
    ._EVAL_18(rsource__EVAL_18),
    ._EVAL_19(rsource__EVAL_19),
    ._EVAL_20(rsource__EVAL_20),
    ._EVAL_21(rsource__EVAL_21),
    ._EVAL_22(rsource__EVAL_22),
    ._EVAL_23(rsource__EVAL_23),
    ._EVAL_24(rsource__EVAL_24),
    ._EVAL_25(rsource__EVAL_25),
    ._EVAL_26(rsource__EVAL_26),
    ._EVAL_27(rsource__EVAL_27),
    ._EVAL_28(rsource__EVAL_28),
    ._EVAL_29(rsource__EVAL_29),
    ._EVAL_30(rsource__EVAL_30),
    ._EVAL_31(rsource__EVAL_31),
    ._EVAL_32(rsource__EVAL_32),
    ._EVAL_33(rsource__EVAL_33),
    ._EVAL_34(rsource__EVAL_34),
    ._EVAL_35(rsource__EVAL_35),
    ._EVAL_36(rsource__EVAL_36),
    ._EVAL_37(rsource__EVAL_37),
    ._EVAL_38(rsource__EVAL_38),
    ._EVAL_39(rsource__EVAL_39),
    ._EVAL_40(rsource__EVAL_40),
    ._EVAL_41(rsource__EVAL_41),
    ._EVAL_42(rsource__EVAL_42),
    ._EVAL_43(rsource__EVAL_43),
    ._EVAL_44(rsource__EVAL_44),
    ._EVAL_45(rsource__EVAL_45),
    ._EVAL_46(rsource__EVAL_46),
    ._EVAL_47(rsource__EVAL_47),
    ._EVAL_48(rsource__EVAL_48),
    ._EVAL_49(rsource__EVAL_49),
    ._EVAL_50(rsource__EVAL_50),
    ._EVAL_51(rsource__EVAL_51),
    ._EVAL_52(rsource__EVAL_52),
    ._EVAL_53(rsource__EVAL_53),
    ._EVAL_54(rsource__EVAL_54),
    ._EVAL_55(rsource__EVAL_55),
    ._EVAL_56(rsource__EVAL_56),
    ._EVAL_57(rsource__EVAL_57),
    ._EVAL_58(rsource__EVAL_58),
    ._EVAL_59(rsource__EVAL_59),
    ._EVAL_60(rsource__EVAL_60),
    ._EVAL_61(rsource__EVAL_61),
    ._EVAL_62(rsource__EVAL_62),
    ._EVAL_63(rsource__EVAL_63),
    ._EVAL_64(rsource__EVAL_64),
    ._EVAL_65(rsource__EVAL_65),
    ._EVAL_66(rsource__EVAL_66),
    ._EVAL_67(rsource__EVAL_67),
    ._EVAL_68(rsource__EVAL_68),
    ._EVAL_69(rsource__EVAL_69),
    ._EVAL_70(rsource__EVAL_70),
    ._EVAL_71(rsource__EVAL_71),
    ._EVAL_72(rsource__EVAL_72),
    ._EVAL_73(rsource__EVAL_73),
    ._EVAL_74(rsource__EVAL_74),
    ._EVAL_75(rsource__EVAL_75),
    ._EVAL_76(rsource__EVAL_76),
    ._EVAL_77(rsource__EVAL_77),
    ._EVAL_78(rsource__EVAL_78),
    ._EVAL_79(rsource__EVAL_79),
    ._EVAL_80(rsource__EVAL_80),
    ._EVAL_81(rsource__EVAL_81),
    ._EVAL_82(rsource__EVAL_82),
    ._EVAL_83(rsource__EVAL_83),
    ._EVAL_84(rsource__EVAL_84),
    ._EVAL_85(rsource__EVAL_85),
    ._EVAL_86(rsource__EVAL_86),
    ._EVAL_87(rsource__EVAL_87),
    ._EVAL_88(rsource__EVAL_88),
    ._EVAL_89(rsource__EVAL_89),
    ._EVAL_90(rsource__EVAL_90),
    ._EVAL_91(rsource__EVAL_91),
    ._EVAL_92(rsource__EVAL_92),
    ._EVAL_93(rsource__EVAL_93),
    ._EVAL_94(rsource__EVAL_94),
    ._EVAL_95(rsource__EVAL_95),
    ._EVAL_96(rsource__EVAL_96),
    ._EVAL_97(rsource__EVAL_97),
    ._EVAL_98(rsource__EVAL_98),
    ._EVAL_99(rsource__EVAL_99),
    ._EVAL_100(rsource__EVAL_100),
    ._EVAL_101(rsource__EVAL_101),
    ._EVAL_102(rsource__EVAL_102),
    ._EVAL_103(rsource__EVAL_103),
    ._EVAL_104(rsource__EVAL_104),
    ._EVAL_105(rsource__EVAL_105),
    ._EVAL_106(rsource__EVAL_106),
    ._EVAL_107(rsource__EVAL_107),
    ._EVAL_108(rsource__EVAL_108)
  );
  SiFive__EVAL_236 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28)
  );
  SiFive__EVAL_287 ptw (
    ._EVAL(ptw__EVAL),
    ._EVAL_0(ptw__EVAL_0),
    ._EVAL_1(ptw__EVAL_1),
    ._EVAL_2(ptw__EVAL_2),
    ._EVAL_3(ptw__EVAL_3),
    ._EVAL_4(ptw__EVAL_4),
    ._EVAL_5(ptw__EVAL_5),
    ._EVAL_6(ptw__EVAL_6),
    ._EVAL_7(ptw__EVAL_7),
    ._EVAL_8(ptw__EVAL_8),
    ._EVAL_9(ptw__EVAL_9),
    ._EVAL_10(ptw__EVAL_10),
    ._EVAL_11(ptw__EVAL_11),
    ._EVAL_12(ptw__EVAL_12),
    ._EVAL_13(ptw__EVAL_13),
    ._EVAL_14(ptw__EVAL_14),
    ._EVAL_15(ptw__EVAL_15),
    ._EVAL_16(ptw__EVAL_16),
    ._EVAL_17(ptw__EVAL_17),
    ._EVAL_18(ptw__EVAL_18),
    ._EVAL_19(ptw__EVAL_19),
    ._EVAL_20(ptw__EVAL_20),
    ._EVAL_21(ptw__EVAL_21),
    ._EVAL_22(ptw__EVAL_22),
    ._EVAL_23(ptw__EVAL_23),
    ._EVAL_24(ptw__EVAL_24),
    ._EVAL_25(ptw__EVAL_25),
    ._EVAL_26(ptw__EVAL_26),
    ._EVAL_27(ptw__EVAL_27),
    ._EVAL_28(ptw__EVAL_28),
    ._EVAL_29(ptw__EVAL_29),
    ._EVAL_30(ptw__EVAL_30),
    ._EVAL_31(ptw__EVAL_31),
    ._EVAL_32(ptw__EVAL_32),
    ._EVAL_33(ptw__EVAL_33),
    ._EVAL_34(ptw__EVAL_34),
    ._EVAL_35(ptw__EVAL_35),
    ._EVAL_36(ptw__EVAL_36),
    ._EVAL_37(ptw__EVAL_37),
    ._EVAL_38(ptw__EVAL_38),
    ._EVAL_39(ptw__EVAL_39),
    ._EVAL_40(ptw__EVAL_40),
    ._EVAL_41(ptw__EVAL_41),
    ._EVAL_42(ptw__EVAL_42),
    ._EVAL_43(ptw__EVAL_43),
    ._EVAL_44(ptw__EVAL_44),
    ._EVAL_45(ptw__EVAL_45),
    ._EVAL_46(ptw__EVAL_46),
    ._EVAL_47(ptw__EVAL_47),
    ._EVAL_48(ptw__EVAL_48),
    ._EVAL_49(ptw__EVAL_49),
    ._EVAL_50(ptw__EVAL_50),
    ._EVAL_51(ptw__EVAL_51),
    ._EVAL_52(ptw__EVAL_52),
    ._EVAL_53(ptw__EVAL_53),
    ._EVAL_54(ptw__EVAL_54),
    ._EVAL_55(ptw__EVAL_55),
    ._EVAL_56(ptw__EVAL_56),
    ._EVAL_57(ptw__EVAL_57),
    ._EVAL_58(ptw__EVAL_58),
    ._EVAL_59(ptw__EVAL_59),
    ._EVAL_60(ptw__EVAL_60),
    ._EVAL_61(ptw__EVAL_61),
    ._EVAL_62(ptw__EVAL_62),
    ._EVAL_63(ptw__EVAL_63),
    ._EVAL_64(ptw__EVAL_64),
    ._EVAL_65(ptw__EVAL_65),
    ._EVAL_66(ptw__EVAL_66),
    ._EVAL_67(ptw__EVAL_67),
    ._EVAL_68(ptw__EVAL_68),
    ._EVAL_69(ptw__EVAL_69),
    ._EVAL_70(ptw__EVAL_70),
    ._EVAL_71(ptw__EVAL_71),
    ._EVAL_72(ptw__EVAL_72),
    ._EVAL_73(ptw__EVAL_73),
    ._EVAL_74(ptw__EVAL_74),
    ._EVAL_75(ptw__EVAL_75),
    ._EVAL_76(ptw__EVAL_76),
    ._EVAL_77(ptw__EVAL_77),
    ._EVAL_78(ptw__EVAL_78),
    ._EVAL_79(ptw__EVAL_79),
    ._EVAL_80(ptw__EVAL_80),
    ._EVAL_81(ptw__EVAL_81),
    ._EVAL_82(ptw__EVAL_82),
    ._EVAL_83(ptw__EVAL_83),
    ._EVAL_84(ptw__EVAL_84),
    ._EVAL_85(ptw__EVAL_85),
    ._EVAL_86(ptw__EVAL_86),
    ._EVAL_87(ptw__EVAL_87),
    ._EVAL_88(ptw__EVAL_88),
    ._EVAL_89(ptw__EVAL_89),
    ._EVAL_90(ptw__EVAL_90),
    ._EVAL_91(ptw__EVAL_91),
    ._EVAL_92(ptw__EVAL_92),
    ._EVAL_93(ptw__EVAL_93),
    ._EVAL_94(ptw__EVAL_94),
    ._EVAL_95(ptw__EVAL_95),
    ._EVAL_96(ptw__EVAL_96),
    ._EVAL_97(ptw__EVAL_97),
    ._EVAL_98(ptw__EVAL_98),
    ._EVAL_99(ptw__EVAL_99),
    ._EVAL_100(ptw__EVAL_100),
    ._EVAL_101(ptw__EVAL_101),
    ._EVAL_102(ptw__EVAL_102),
    ._EVAL_103(ptw__EVAL_103),
    ._EVAL_104(ptw__EVAL_104),
    ._EVAL_105(ptw__EVAL_105),
    ._EVAL_106(ptw__EVAL_106),
    ._EVAL_107(ptw__EVAL_107),
    ._EVAL_108(ptw__EVAL_108),
    ._EVAL_109(ptw__EVAL_109),
    ._EVAL_110(ptw__EVAL_110),
    ._EVAL_111(ptw__EVAL_111),
    ._EVAL_112(ptw__EVAL_112),
    ._EVAL_113(ptw__EVAL_113),
    ._EVAL_114(ptw__EVAL_114),
    ._EVAL_115(ptw__EVAL_115),
    ._EVAL_116(ptw__EVAL_116),
    ._EVAL_117(ptw__EVAL_117),
    ._EVAL_118(ptw__EVAL_118),
    ._EVAL_119(ptw__EVAL_119),
    ._EVAL_120(ptw__EVAL_120),
    ._EVAL_121(ptw__EVAL_121),
    ._EVAL_122(ptw__EVAL_122),
    ._EVAL_123(ptw__EVAL_123),
    ._EVAL_124(ptw__EVAL_124),
    ._EVAL_125(ptw__EVAL_125),
    ._EVAL_126(ptw__EVAL_126),
    ._EVAL_127(ptw__EVAL_127),
    ._EVAL_128(ptw__EVAL_128),
    ._EVAL_129(ptw__EVAL_129),
    ._EVAL_130(ptw__EVAL_130),
    ._EVAL_131(ptw__EVAL_131),
    ._EVAL_132(ptw__EVAL_132),
    ._EVAL_133(ptw__EVAL_133),
    ._EVAL_134(ptw__EVAL_134),
    ._EVAL_135(ptw__EVAL_135),
    ._EVAL_136(ptw__EVAL_136),
    ._EVAL_137(ptw__EVAL_137),
    ._EVAL_138(ptw__EVAL_138),
    ._EVAL_139(ptw__EVAL_139),
    ._EVAL_140(ptw__EVAL_140),
    ._EVAL_141(ptw__EVAL_141),
    ._EVAL_142(ptw__EVAL_142),
    ._EVAL_143(ptw__EVAL_143),
    ._EVAL_144(ptw__EVAL_144),
    ._EVAL_145(ptw__EVAL_145),
    ._EVAL_146(ptw__EVAL_146),
    ._EVAL_147(ptw__EVAL_147),
    ._EVAL_148(ptw__EVAL_148),
    ._EVAL_149(ptw__EVAL_149),
    ._EVAL_150(ptw__EVAL_150),
    ._EVAL_151(ptw__EVAL_151),
    ._EVAL_152(ptw__EVAL_152),
    ._EVAL_153(ptw__EVAL_153),
    ._EVAL_154(ptw__EVAL_154),
    ._EVAL_155(ptw__EVAL_155),
    ._EVAL_156(ptw__EVAL_156),
    ._EVAL_157(ptw__EVAL_157),
    ._EVAL_158(ptw__EVAL_158),
    ._EVAL_159(ptw__EVAL_159),
    ._EVAL_160(ptw__EVAL_160),
    ._EVAL_161(ptw__EVAL_161),
    ._EVAL_162(ptw__EVAL_162),
    ._EVAL_163(ptw__EVAL_163),
    ._EVAL_164(ptw__EVAL_164),
    ._EVAL_165(ptw__EVAL_165),
    ._EVAL_166(ptw__EVAL_166),
    ._EVAL_167(ptw__EVAL_167),
    ._EVAL_168(ptw__EVAL_168),
    ._EVAL_169(ptw__EVAL_169),
    ._EVAL_170(ptw__EVAL_170),
    ._EVAL_171(ptw__EVAL_171),
    ._EVAL_172(ptw__EVAL_172),
    ._EVAL_173(ptw__EVAL_173),
    ._EVAL_174(ptw__EVAL_174),
    ._EVAL_175(ptw__EVAL_175),
    ._EVAL_176(ptw__EVAL_176),
    ._EVAL_177(ptw__EVAL_177),
    ._EVAL_178(ptw__EVAL_178),
    ._EVAL_179(ptw__EVAL_179)
  );
  SiFive__EVAL_234 frontend (
    ._EVAL(frontend__EVAL),
    ._EVAL_0(frontend__EVAL_0),
    ._EVAL_1(frontend__EVAL_1),
    ._EVAL_2(frontend__EVAL_2),
    ._EVAL_3(frontend__EVAL_3),
    ._EVAL_4(frontend__EVAL_4),
    ._EVAL_5(frontend__EVAL_5),
    ._EVAL_6(frontend__EVAL_6),
    ._EVAL_7(frontend__EVAL_7),
    ._EVAL_8(frontend__EVAL_8),
    ._EVAL_9(frontend__EVAL_9),
    ._EVAL_10(frontend__EVAL_10),
    ._EVAL_11(frontend__EVAL_11),
    ._EVAL_12(frontend__EVAL_12),
    ._EVAL_13(frontend__EVAL_13),
    ._EVAL_14(frontend__EVAL_14),
    ._EVAL_15(frontend__EVAL_15),
    ._EVAL_16(frontend__EVAL_16),
    ._EVAL_17(frontend__EVAL_17),
    ._EVAL_18(frontend__EVAL_18),
    ._EVAL_19(frontend__EVAL_19),
    ._EVAL_20(frontend__EVAL_20),
    ._EVAL_21(frontend__EVAL_21),
    ._EVAL_22(frontend__EVAL_22),
    ._EVAL_23(frontend__EVAL_23),
    ._EVAL_24(frontend__EVAL_24),
    ._EVAL_25(frontend__EVAL_25),
    ._EVAL_26(frontend__EVAL_26),
    ._EVAL_27(frontend__EVAL_27),
    ._EVAL_28(frontend__EVAL_28),
    ._EVAL_29(frontend__EVAL_29),
    ._EVAL_30(frontend__EVAL_30),
    ._EVAL_31(frontend__EVAL_31),
    ._EVAL_32(frontend__EVAL_32),
    ._EVAL_33(frontend__EVAL_33),
    ._EVAL_34(frontend__EVAL_34),
    ._EVAL_35(frontend__EVAL_35),
    ._EVAL_36(frontend__EVAL_36),
    ._EVAL_37(frontend__EVAL_37),
    ._EVAL_38(frontend__EVAL_38),
    ._EVAL_39(frontend__EVAL_39),
    ._EVAL_40(frontend__EVAL_40),
    ._EVAL_41(frontend__EVAL_41),
    ._EVAL_42(frontend__EVAL_42),
    ._EVAL_43(frontend__EVAL_43),
    ._EVAL_44(frontend__EVAL_44),
    ._EVAL_45(frontend__EVAL_45),
    ._EVAL_46(frontend__EVAL_46),
    ._EVAL_47(frontend__EVAL_47),
    ._EVAL_48(frontend__EVAL_48),
    ._EVAL_49(frontend__EVAL_49),
    ._EVAL_50(frontend__EVAL_50),
    ._EVAL_51(frontend__EVAL_51),
    ._EVAL_52(frontend__EVAL_52),
    ._EVAL_53(frontend__EVAL_53),
    ._EVAL_54(frontend__EVAL_54),
    ._EVAL_55(frontend__EVAL_55),
    ._EVAL_56(frontend__EVAL_56),
    ._EVAL_57(frontend__EVAL_57),
    ._EVAL_58(frontend__EVAL_58),
    ._EVAL_59(frontend__EVAL_59),
    ._EVAL_60(frontend__EVAL_60),
    ._EVAL_61(frontend__EVAL_61),
    ._EVAL_62(frontend__EVAL_62),
    ._EVAL_63(frontend__EVAL_63),
    ._EVAL_64(frontend__EVAL_64),
    ._EVAL_65(frontend__EVAL_65),
    ._EVAL_66(frontend__EVAL_66),
    ._EVAL_67(frontend__EVAL_67),
    ._EVAL_68(frontend__EVAL_68),
    ._EVAL_69(frontend__EVAL_69),
    ._EVAL_70(frontend__EVAL_70),
    ._EVAL_71(frontend__EVAL_71),
    ._EVAL_72(frontend__EVAL_72),
    ._EVAL_73(frontend__EVAL_73),
    ._EVAL_74(frontend__EVAL_74),
    ._EVAL_75(frontend__EVAL_75),
    ._EVAL_76(frontend__EVAL_76),
    ._EVAL_77(frontend__EVAL_77),
    ._EVAL_78(frontend__EVAL_78),
    ._EVAL_79(frontend__EVAL_79),
    ._EVAL_80(frontend__EVAL_80),
    ._EVAL_81(frontend__EVAL_81),
    ._EVAL_82(frontend__EVAL_82),
    ._EVAL_83(frontend__EVAL_83),
    ._EVAL_84(frontend__EVAL_84),
    ._EVAL_85(frontend__EVAL_85),
    ._EVAL_86(frontend__EVAL_86),
    ._EVAL_87(frontend__EVAL_87),
    ._EVAL_88(frontend__EVAL_88),
    ._EVAL_89(frontend__EVAL_89),
    ._EVAL_90(frontend__EVAL_90),
    ._EVAL_91(frontend__EVAL_91),
    ._EVAL_92(frontend__EVAL_92),
    ._EVAL_93(frontend__EVAL_93),
    ._EVAL_94(frontend__EVAL_94),
    ._EVAL_95(frontend__EVAL_95),
    ._EVAL_96(frontend__EVAL_96),
    ._EVAL_97(frontend__EVAL_97),
    ._EVAL_98(frontend__EVAL_98),
    ._EVAL_99(frontend__EVAL_99),
    ._EVAL_100(frontend__EVAL_100),
    ._EVAL_101(frontend__EVAL_101),
    ._EVAL_102(frontend__EVAL_102),
    ._EVAL_103(frontend__EVAL_103),
    ._EVAL_104(frontend__EVAL_104),
    ._EVAL_105(frontend__EVAL_105),
    ._EVAL_106(frontend__EVAL_106),
    ._EVAL_107(frontend__EVAL_107),
    ._EVAL_108(frontend__EVAL_108),
    ._EVAL_109(frontend__EVAL_109),
    ._EVAL_110(frontend__EVAL_110),
    ._EVAL_111(frontend__EVAL_111),
    ._EVAL_112(frontend__EVAL_112),
    ._EVAL_113(frontend__EVAL_113),
    ._EVAL_114(frontend__EVAL_114),
    ._EVAL_115(frontend__EVAL_115),
    ._EVAL_116(frontend__EVAL_116),
    ._EVAL_117(frontend__EVAL_117),
    ._EVAL_118(frontend__EVAL_118),
    ._EVAL_119(frontend__EVAL_119),
    ._EVAL_120(frontend__EVAL_120),
    ._EVAL_121(frontend__EVAL_121),
    ._EVAL_122(frontend__EVAL_122),
    ._EVAL_123(frontend__EVAL_123),
    ._EVAL_124(frontend__EVAL_124),
    ._EVAL_125(frontend__EVAL_125),
    ._EVAL_126(frontend__EVAL_126),
    ._EVAL_127(frontend__EVAL_127),
    ._EVAL_128(frontend__EVAL_128),
    ._EVAL_129(frontend__EVAL_129),
    ._EVAL_130(frontend__EVAL_130),
    ._EVAL_131(frontend__EVAL_131),
    ._EVAL_132(frontend__EVAL_132),
    ._EVAL_133(frontend__EVAL_133),
    ._EVAL_134(frontend__EVAL_134),
    ._EVAL_135(frontend__EVAL_135),
    ._EVAL_136(frontend__EVAL_136),
    ._EVAL_137(frontend__EVAL_137),
    ._EVAL_138(frontend__EVAL_138),
    ._EVAL_139(frontend__EVAL_139),
    ._EVAL_140(frontend__EVAL_140),
    ._EVAL_141(frontend__EVAL_141),
    ._EVAL_142(frontend__EVAL_142)
  );
  SiFive__EVAL_277 rsink (
    ._EVAL(rsink__EVAL),
    ._EVAL_0(rsink__EVAL_0),
    ._EVAL_1(rsink__EVAL_1),
    ._EVAL_2(rsink__EVAL_2),
    ._EVAL_3(rsink__EVAL_3),
    ._EVAL_4(rsink__EVAL_4),
    ._EVAL_5(rsink__EVAL_5),
    ._EVAL_6(rsink__EVAL_6),
    ._EVAL_7(rsink__EVAL_7),
    ._EVAL_8(rsink__EVAL_8),
    ._EVAL_9(rsink__EVAL_9),
    ._EVAL_10(rsink__EVAL_10),
    ._EVAL_11(rsink__EVAL_11),
    ._EVAL_12(rsink__EVAL_12),
    ._EVAL_13(rsink__EVAL_13),
    ._EVAL_14(rsink__EVAL_14),
    ._EVAL_15(rsink__EVAL_15),
    ._EVAL_16(rsink__EVAL_16),
    ._EVAL_17(rsink__EVAL_17),
    ._EVAL_18(rsink__EVAL_18),
    ._EVAL_19(rsink__EVAL_19),
    ._EVAL_20(rsink__EVAL_20),
    ._EVAL_21(rsink__EVAL_21),
    ._EVAL_22(rsink__EVAL_22),
    ._EVAL_23(rsink__EVAL_23),
    ._EVAL_24(rsink__EVAL_24),
    ._EVAL_25(rsink__EVAL_25),
    ._EVAL_26(rsink__EVAL_26),
    ._EVAL_27(rsink__EVAL_27),
    ._EVAL_28(rsink__EVAL_28),
    ._EVAL_29(rsink__EVAL_29),
    ._EVAL_30(rsink__EVAL_30),
    ._EVAL_31(rsink__EVAL_31),
    ._EVAL_32(rsink__EVAL_32),
    ._EVAL_33(rsink__EVAL_33),
    ._EVAL_34(rsink__EVAL_34),
    ._EVAL_35(rsink__EVAL_35),
    ._EVAL_36(rsink__EVAL_36),
    ._EVAL_37(rsink__EVAL_37),
    ._EVAL_38(rsink__EVAL_38),
    ._EVAL_39(rsink__EVAL_39),
    ._EVAL_40(rsink__EVAL_40),
    ._EVAL_41(rsink__EVAL_41),
    ._EVAL_42(rsink__EVAL_42),
    ._EVAL_43(rsink__EVAL_43),
    ._EVAL_44(rsink__EVAL_44),
    ._EVAL_45(rsink__EVAL_45),
    ._EVAL_46(rsink__EVAL_46),
    ._EVAL_47(rsink__EVAL_47),
    ._EVAL_48(rsink__EVAL_48),
    ._EVAL_49(rsink__EVAL_49),
    ._EVAL_50(rsink__EVAL_50),
    ._EVAL_51(rsink__EVAL_51),
    ._EVAL_52(rsink__EVAL_52),
    ._EVAL_53(rsink__EVAL_53),
    ._EVAL_54(rsink__EVAL_54),
    ._EVAL_55(rsink__EVAL_55),
    ._EVAL_56(rsink__EVAL_56),
    ._EVAL_57(rsink__EVAL_57),
    ._EVAL_58(rsink__EVAL_58),
    ._EVAL_59(rsink__EVAL_59),
    ._EVAL_60(rsink__EVAL_60)
  );
  SiFive__EVAL_246 dlsXbar (
    ._EVAL(dlsXbar__EVAL),
    ._EVAL_0(dlsXbar__EVAL_0),
    ._EVAL_1(dlsXbar__EVAL_1),
    ._EVAL_2(dlsXbar__EVAL_2),
    ._EVAL_3(dlsXbar__EVAL_3),
    ._EVAL_4(dlsXbar__EVAL_4),
    ._EVAL_5(dlsXbar__EVAL_5),
    ._EVAL_6(dlsXbar__EVAL_6),
    ._EVAL_7(dlsXbar__EVAL_7),
    ._EVAL_8(dlsXbar__EVAL_8),
    ._EVAL_9(dlsXbar__EVAL_9),
    ._EVAL_10(dlsXbar__EVAL_10),
    ._EVAL_11(dlsXbar__EVAL_11),
    ._EVAL_12(dlsXbar__EVAL_12),
    ._EVAL_13(dlsXbar__EVAL_13),
    ._EVAL_14(dlsXbar__EVAL_14),
    ._EVAL_15(dlsXbar__EVAL_15),
    ._EVAL_16(dlsXbar__EVAL_16),
    ._EVAL_17(dlsXbar__EVAL_17),
    ._EVAL_18(dlsXbar__EVAL_18),
    ._EVAL_19(dlsXbar__EVAL_19),
    ._EVAL_20(dlsXbar__EVAL_20),
    ._EVAL_21(dlsXbar__EVAL_21),
    ._EVAL_22(dlsXbar__EVAL_22),
    ._EVAL_23(dlsXbar__EVAL_23),
    ._EVAL_24(dlsXbar__EVAL_24),
    ._EVAL_25(dlsXbar__EVAL_25),
    ._EVAL_26(dlsXbar__EVAL_26),
    ._EVAL_27(dlsXbar__EVAL_27),
    ._EVAL_28(dlsXbar__EVAL_28),
    ._EVAL_29(dlsXbar__EVAL_29),
    ._EVAL_30(dlsXbar__EVAL_30),
    ._EVAL_31(dlsXbar__EVAL_31),
    ._EVAL_32(dlsXbar__EVAL_32),
    ._EVAL_33(dlsXbar__EVAL_33),
    ._EVAL_34(dlsXbar__EVAL_34),
    ._EVAL_35(dlsXbar__EVAL_35),
    ._EVAL_36(dlsXbar__EVAL_36),
    ._EVAL_37(dlsXbar__EVAL_37),
    ._EVAL_38(dlsXbar__EVAL_38),
    ._EVAL_39(dlsXbar__EVAL_39),
    ._EVAL_40(dlsXbar__EVAL_40),
    ._EVAL_41(dlsXbar__EVAL_41),
    ._EVAL_42(dlsXbar__EVAL_42),
    ._EVAL_43(dlsXbar__EVAL_43),
    ._EVAL_44(dlsXbar__EVAL_44),
    ._EVAL_45(dlsXbar__EVAL_45),
    ._EVAL_46(dlsXbar__EVAL_46),
    ._EVAL_47(dlsXbar__EVAL_47),
    ._EVAL_48(dlsXbar__EVAL_48)
  );
  assign core__EVAL_196 = dcacheArb__EVAL_89;
  assign buffer_1__EVAL_22 = dlsXbar__EVAL_39;
  assign InstructionQueue__EVAL_15 = FormMicroOps__EVAL_121;
  assign filter__EVAL_53 = tlMasterXbar__EVAL_24;
  assign rsource__EVAL_62 = buffer_2__EVAL_22;
  assign buffer_2__EVAL_8 = tlMasterXbar__EVAL_48;
  assign intsink_2__EVAL_0 = _EVAL_24;
  assign core__EVAL_81 = dcacheArb__EVAL_68;
  assign filter__EVAL_38 = coreXbar__EVAL_51;
  assign dcache__EVAL_150 = ptw__EVAL_160;
  assign buffer__EVAL = tlMasterXbar__EVAL_73;
  assign FormMicroOps__EVAL_154 = core__EVAL_219;
  assign ptw__EVAL_115 = core__EVAL_181;
  assign rsource__EVAL_102 = _EVAL_0;
  assign frontend__EVAL_20 = core__EVAL_75;
  assign frontend__EVAL_80 = core__EVAL_229;
  assign FormMicroOps__EVAL_143 = frontend__EVAL_111;
  assign rsink__EVAL_21 = _EVAL_32;
  assign dls__EVAL_12 = fragmenter_1__EVAL_30;
  assign dcache__EVAL_28 = ptw__EVAL_10;
  assign dcache__EVAL_39 = ptw__EVAL_95;
  assign tlMasterXbar__EVAL_9 = filter__EVAL_23;
  assign widget__EVAL_12 = _EVAL_32;
  assign frontend__EVAL_40 = ptw__EVAL_91;
  assign frontend__EVAL_134 = ptw__EVAL_176;
  assign frontend__EVAL_138 = core__EVAL_244;
  assign coreXbar__EVAL_1 = dcache__EVAL_121;
  assign core__EVAL_23 = InstructionQueue__EVAL_152;
  assign filter__EVAL_11 = tlMasterXbar__EVAL_0;
  assign frontend__EVAL_47 = ptw__EVAL_32;
  assign core__EVAL_249 = dcacheArb__EVAL_31;
  assign core__EVAL_268 = InstructionQueue__EVAL_173;
  assign dlsXbar__EVAL_16 = widget_1__EVAL_22;
  assign dcache__EVAL_104 = dcacheArb__EVAL_78;
  assign frontend__EVAL_34 = core__EVAL_218;
  assign filter__EVAL_61 = coreXbar__EVAL_46;
  assign FormMicroOps__EVAL_53 = core__EVAL_144;
  assign dcache__EVAL_141 = ptw__EVAL_9;
  assign frontend__EVAL_94 = core__EVAL_238;
  assign rsource__EVAL_108 = _EVAL_102;
  assign dcache__EVAL_11 = ptw__EVAL_51;
  assign _EVAL_99 = rsource__EVAL_63;
  assign ptw__EVAL_177 = core__EVAL_72;
  assign ptw__EVAL_72 = core__EVAL_67;
  assign core__EVAL_165 = InstructionQueue__EVAL_132;
  assign widget__EVAL_11 = tlSlaveXbar__EVAL_46;
  assign fragmenter_1__EVAL_20 = dls__EVAL_13;
  assign frontend__EVAL_46 = core__EVAL_258;
  assign coreXbar__EVAL_70 = widget_1__EVAL_24;
  assign buffer_1__EVAL_20 = dlsXbar__EVAL_29;
  assign ptw__EVAL_165 = core__EVAL_11;
  assign rsource__EVAL_67 = buffer_2__EVAL_33;
  assign buffer_2__EVAL_40 = rsource__EVAL_49;
  assign tlSlaveXbar__EVAL_23 = widget__EVAL;
  assign rsink__EVAL_35 = _EVAL_48;
  assign core__EVAL_90 = InstructionQueue__EVAL_43;
  assign frontend__EVAL_136 = ptw__EVAL_85;
  assign FormMicroOps__EVAL_73 = frontend__EVAL_91;
  assign dcacheArb__EVAL_72 = core__EVAL_38;
  assign frontend__EVAL_123 = ptw__EVAL_46;
  assign dlsXbar__EVAL_14 = buffer_1__EVAL_5;
  assign core__EVAL_168 = InstructionQueue__EVAL_159;
  assign core__EVAL_224 = InstructionQueue__EVAL_21;
  assign coreXbar__EVAL_20 = dcache__EVAL_70;
  assign core__EVAL_172 = InstructionQueue__EVAL_106;
  assign dlsXbar__EVAL_5 = buffer_1__EVAL_25;
  assign frontend__EVAL_41 = ptw__EVAL_143;
  assign frontend__EVAL_119 = ptw__EVAL_163;
  assign InstructionQueue__EVAL_39 = FormMicroOps__EVAL_93;
  assign frontend__EVAL_116 = core__EVAL_13;
  assign frontend__EVAL_122 = buffer__EVAL_0;
  assign tlMasterXbar__EVAL_60 = buffer__EVAL_14;
  assign buffer__EVAL_13 = tlMasterXbar__EVAL_69;
  assign tlSlaveXbar__EVAL_42 = widget__EVAL_10;
  assign filter__EVAL_51 = tlMasterXbar__EVAL_8;
  assign core__EVAL_51 = InstructionQueue__EVAL_24;
  assign dcache__EVAL_62 = ptw__EVAL_113;
  assign FormMicroOps__EVAL_126 = core__EVAL_166;
  assign core__EVAL_40 = InstructionQueue__EVAL_17;
  assign core__EVAL_278 = InstructionQueue__EVAL_38;
  assign FormMicroOps__EVAL_67 = core__EVAL_70;
  assign dcache__EVAL_102 = ptw__EVAL_17;
  assign core__EVAL_35 = InstructionQueue__EVAL_67;
  assign coreXbar__EVAL_67 = filter__EVAL_62;
  assign dlsXbar__EVAL_35 = _EVAL_32;
  assign FormMicroOps__EVAL_89 = core__EVAL_101;
  assign fragmenter_1__EVAL_27 = buffer_1__EVAL;
  assign _EVAL_88 = rsource__EVAL_19;
  assign tlMasterXbar__EVAL_6 = filter__EVAL_30;
  assign core__EVAL_142 = dcacheArb__EVAL_86;
  assign buffer_1__EVAL_19 = dlsXbar__EVAL_23;
  assign buffer_2__EVAL_16 = tlMasterXbar__EVAL_54;
  assign buffer_2__EVAL_44 = rsource__EVAL_10;
  assign tlMasterXbar__EVAL_3 = filter__EVAL_31;
  assign FormMicroOps__EVAL_98 = core__EVAL_241;
  assign core__EVAL_208 = InstructionQueue__EVAL_30;
  assign core__EVAL_55 = InstructionQueue__EVAL_56;
  assign _EVAL_66 = rsource__EVAL_80;
  assign _EVAL_93 = rsource__EVAL_20;
  assign rsource__EVAL_78 = _EVAL_31;
  assign buffer_3__EVAL_12 = tlSlaveXbar__EVAL_24;
  assign frontend__EVAL_98 = ptw__EVAL_55;
  assign InstructionQueue__EVAL_99 = FormMicroOps__EVAL_159;
  assign rsource__EVAL_86 = _EVAL_30;
  assign dcacheArb__EVAL_88 = dcache__EVAL_43;
  assign dcache__EVAL_148 = dcacheArb__EVAL_55;
  assign buffer__EVAL_5 = tlMasterXbar__EVAL_21;
  assign FormMicroOps__EVAL_104 = core__EVAL_152;
  assign tlMasterXbar__EVAL_14 = filter__EVAL_25;
  assign dlsXbar__EVAL_24 = widget_1__EVAL_31;
  assign InstructionQueue__EVAL_92 = FormMicroOps__EVAL_10;
  assign filter__EVAL_14 = tlMasterXbar__EVAL_33;
  assign core__EVAL_110 = dcacheArb__EVAL_32;
  assign coreXbar__EVAL_54 = widget_1__EVAL_28;
  assign rsource__EVAL_107 = _EVAL_68;
  assign frontend__EVAL_103 = buffer__EVAL_8;
  assign _EVAL_3 = rsource__EVAL_6;
  assign buffer_1__EVAL_14 = dlsXbar__EVAL_47;
  assign tlMasterXbar__EVAL_61 = filter__EVAL_19;
  assign core__EVAL_246 = dcacheArb__EVAL_6;
  assign dcache__EVAL_133 = dcacheArb__EVAL_81;
  assign frontend__EVAL_95 = ptw__EVAL_154;
  assign core__EVAL_16 = InstructionQueue__EVAL_136;
  assign ptw__EVAL_13 = core__EVAL_88;
  assign fragmenter__EVAL_7 = frontend__EVAL_120;
  assign core__EVAL_122 = dcacheArb__EVAL_58;
  assign buffer_1__EVAL_17 = fragmenter_1__EVAL_5;
  assign filter__EVAL_71 = coreXbar__EVAL_31;
  assign InstructionQueue__EVAL_105 = FormMicroOps__EVAL_99;
  assign core__EVAL_127 = _EVAL_67;
  assign fragmenter_1__EVAL_2 = _EVAL_100;
  assign coreXbar__EVAL = dcache__EVAL_59;
  assign frontend__EVAL_21 = ptw__EVAL_78;
  assign _EVAL_37 = rsource__EVAL_36;
  assign fragmenter__EVAL_12 = widget__EVAL_7;
  assign frontend__EVAL_18 = core__EVAL_93;
  assign ptw__EVAL_169 = core__EVAL_44;
  assign widget_1__EVAL_14 = dlsXbar__EVAL_36;
  assign widget_1__EVAL_16 = coreXbar__EVAL_37;
  assign widget_1__EVAL_19 = coreXbar__EVAL_55;
  assign core__EVAL_188 = InstructionQueue__EVAL_26;
  assign ptw__EVAL_119 = core__EVAL_256;
  assign rsource__EVAL_54 = _EVAL_94;
  assign _EVAL_77 = rsink__EVAL_30;
  assign ptw__EVAL_98 = core__EVAL_89;
  assign InstructionQueue__EVAL_42 = FormMicroOps__EVAL_113;
  assign widget__EVAL_24 = tlSlaveXbar__EVAL_47;
  assign buffer_2__EVAL_35 = tlMasterXbar__EVAL_7;
  assign frontend__EVAL_93 = ptw__EVAL_122;
  assign dcache__EVAL_60 = ptw__EVAL_106;
  assign FormMicroOps__EVAL_51 = _EVAL_100;
  assign tlMasterXbar__EVAL_53 = filter__EVAL_24;
  assign dlsXbar__EVAL_15 = buffer_1__EVAL_23;
  assign tlSlaveXbar__EVAL_11 = buffer_3__EVAL_0;
  assign rsink__EVAL_22 = _EVAL_90;
  assign coreXbar__EVAL_8 = filter__EVAL_10;
  assign dcacheArb__EVAL_14 = dcache__EVAL_111;
  assign _EVAL_11 = rsource__EVAL_92;
  assign _EVAL_27 = rsource__EVAL_0;
  assign buffer_3__EVAL_28 = tlSlaveXbar__EVAL_13;
  assign fragmenter_1__EVAL_28 = dls__EVAL_7;
  assign frontend__EVAL_140 = ptw__EVAL_131;
  assign buffer_2__EVAL_18 = tlMasterXbar__EVAL_57;
  assign dcacheArb__EVAL_54 = dcache__EVAL_91;
  assign rsource__EVAL_27 = _EVAL_2;
  assign coreXbar__EVAL_48 = filter__EVAL_65;
  assign InstructionQueue__EVAL_46 = FormMicroOps__EVAL_78;
  assign coreXbar__EVAL_83 = filter__EVAL_34;
  assign FormMicroOps__EVAL_42 = frontend__EVAL_127;
  assign dcacheArb__EVAL_9 = dcache__EVAL_108;
  assign FormMicroOps__EVAL_64 = core__EVAL_210;
  assign filter__EVAL_72 = coreXbar__EVAL_30;
  assign rsource__EVAL_52 = _EVAL_14;
  assign core__EVAL_251 = InstructionQueue__EVAL_65;
  assign FormMicroOps__EVAL_52 = frontend__EVAL_135;
  assign dcache__EVAL_54 = dcacheArb__EVAL_53;
  assign InstructionQueue__EVAL_139 = FormMicroOps__EVAL_138;
  assign core__EVAL_198 = InstructionQueue__EVAL_59;
  assign frontend__EVAL_97 = buffer__EVAL_15;
  assign dcache__EVAL_83 = ptw__EVAL_128;
  assign ptw__EVAL_159 = core__EVAL_10;
  assign FormMicroOps__EVAL_44 = core__EVAL_162;
  assign rsink__EVAL_39 = _EVAL_28;
  assign FormMicroOps__EVAL_24 = core__EVAL_227;
  assign fragmenter_1__EVAL_9 = buffer_1__EVAL_12;
  assign FormMicroOps__EVAL_1 = frontend__EVAL_1;
  assign dcacheArb__EVAL_30 = dcache__EVAL_64;
  assign frontend__EVAL_77 = core__EVAL_54;
  assign core__EVAL_206 = InstructionQueue__EVAL_134;
  assign dlsXbar__EVAL_42 = tlSlaveXbar__EVAL_40;
  assign core__EVAL_159 = dcacheArb__EVAL_67;
  assign InstructionQueue__EVAL_143 = FormMicroOps__EVAL_58;
  assign frontend__EVAL_115 = ptw__EVAL_25;
  assign _EVAL_57 = rsource__EVAL_48;
  assign frontend__EVAL_128 = ptw__EVAL_103;
  assign _EVAL_96 = rsource__EVAL_37;
  assign coreXbar__EVAL_2 = dcache__EVAL_100;
  assign dlsXbar__EVAL_7 = tlSlaveXbar__EVAL_34;
  assign dlsXbar__EVAL_26 = widget_1__EVAL_27;
  assign core__EVAL_107 = dcacheArb__EVAL_33;
  assign dcache__EVAL_67 = ptw__EVAL_89;
  assign rsource__EVAL_84 = _EVAL_115;
  assign buffer_3__EVAL_14 = tlSlaveXbar__EVAL_22;
  assign dlsXbar__EVAL_31 = buffer_1__EVAL_24;
  assign buffer_1__EVAL_8 = _EVAL_32;
  assign FormMicroOps__EVAL_39 = core__EVAL_28;
  assign core__EVAL_215 = dcacheArb__EVAL_51;
  assign core__EVAL_232 = InstructionQueue__EVAL_83;
  assign widget_1__EVAL_9 = coreXbar__EVAL_57;
  assign intsink__EVAL_1 = _EVAL_80;
  assign tlSlaveXbar__EVAL_50 = widget__EVAL_28;
  assign _EVAL_18 = rsource__EVAL_64;
  assign _EVAL_15 = rsource__EVAL_58;
  assign dcacheArb__EVAL_65 = core__EVAL_5;
  assign dcache__EVAL_77 = 4'h0;
  assign core__EVAL_102 = InstructionQueue__EVAL_180;
  assign core__EVAL_176 = InstructionQueue__EVAL_70;
  assign ptw__EVAL_179 = core__EVAL_77;
  assign core__EVAL_15 = dcacheArb__EVAL_79;
  assign rsink__EVAL_15 = buffer_3__EVAL_1;
  assign InstructionQueue__EVAL_135 = FormMicroOps__EVAL_87;
  assign tlMasterXbar__EVAL_46 = buffer_2__EVAL_57;
  assign rsink__EVAL_13 = _EVAL_8;
  assign core__EVAL_267 = _EVAL_100;
  assign buffer_2__EVAL_37 = _EVAL_100;
  assign dcache__EVAL_71 = dcacheArb__EVAL_13;
  assign rsource__EVAL_26 = buffer_2__EVAL_69;
  assign tlSlaveXbar__EVAL_31 = buffer_3__EVAL_2;
  assign dlsXbar__EVAL_20 = widget_1__EVAL_29;
  assign _EVAL_1 = rsink__EVAL_4;
  assign _EVAL_10 = rsource__EVAL_57;
  assign rsink__EVAL_47 = buffer_3__EVAL_13;
  assign dcacheArb__EVAL_35 = dcache__EVAL_17;
  assign tlMasterXbar__EVAL_74 = filter__EVAL_29;
  assign dcache__EVAL_10 = coreXbar__EVAL_60;
  assign dcacheArb__EVAL_37 = dcache__EVAL_47;
  assign InstructionQueue__EVAL_120 = FormMicroOps__EVAL_11;
  assign core__EVAL_138 = InstructionQueue__EVAL_146;
  assign dcache__EVAL_19 = ptw__EVAL_102;
  assign _EVAL_29 = rsource__EVAL_8;
  assign _EVAL_65 = rsink__EVAL_17;
  assign buffer_2__EVAL_1 = rsource__EVAL_72;
  assign ptw__EVAL_38 = core__EVAL_178;
  assign rsource__EVAL_69 = buffer_2__EVAL_13;
  assign InstructionQueue__EVAL_122 = FormMicroOps__EVAL_16;
  assign dlsXbar__EVAL_19 = tlSlaveXbar__EVAL_21;
  assign dcache__EVAL_49 = coreXbar__EVAL_61;
  assign InstructionQueue__EVAL_35 = FormMicroOps__EVAL_140;
  assign frontend__EVAL_36 = core__EVAL_114;
  assign _EVAL_46 = rsource__EVAL_85;
  assign _EVAL_79 = rsource__EVAL_2;
  assign dlsXbar__EVAL_44 = tlSlaveXbar__EVAL_37;
  assign rsink__EVAL_43 = _EVAL_104;
  assign filter__EVAL_35 = coreXbar__EVAL_44;
  assign rsource__EVAL_96 = buffer_2__EVAL_39;
  assign dcache__EVAL_37 = dcacheArb__EVAL_87;
  assign coreXbar__EVAL_49 = dcache__EVAL_30;
  assign fragmenter_1__EVAL_18 = buffer_1__EVAL_15;
  assign ptw__EVAL_16 = core__EVAL_48;
  assign InstructionQueue__EVAL_149 = FormMicroOps__EVAL_148;
  assign filter__EVAL_33 = tlMasterXbar__EVAL_12;
  assign tlMasterXbar__EVAL_19 = filter__EVAL_50;
  assign core__EVAL_97 = InstructionQueue__EVAL_98;
  assign dls__EVAL_6 = fragmenter_1__EVAL_8;
  assign core__EVAL_154 = InstructionQueue__EVAL_27;
  assign fragmenter_1__EVAL_0 = buffer_1__EVAL_30;
  assign buffer_1__EVAL_28 = fragmenter_1__EVAL_3;
  assign dcache__EVAL_29 = ptw__EVAL_47;
  assign core__EVAL_203 = dcacheArb__EVAL_84;
  assign dlsXbar__EVAL_8 = tlSlaveXbar__EVAL_19;
  assign ptw__EVAL_7 = core__EVAL_230;
  assign ptw__EVAL_77 = core__EVAL_130;
  assign ptw__EVAL_52 = core__EVAL_125;
  assign buffer_2__EVAL_60 = tlMasterXbar__EVAL_32;
  assign core__EVAL_59 = InstructionQueue__EVAL_185;
  assign dcacheArb__EVAL_39 = core__EVAL_50;
  assign filter__EVAL_44 = tlMasterXbar__EVAL_72;
  assign FormMicroOps__EVAL_132 = core__EVAL_157;
  assign rsink__EVAL_41 = _EVAL_63;
  assign frontend__EVAL_88 = ptw__EVAL_71;
  assign dcache__EVAL_95 = ptw__EVAL_173;
  assign core__EVAL_119 = InstructionQueue__EVAL_170;
  assign ptw__EVAL_84 = core__EVAL_37;
  assign rsource__EVAL_4 = buffer_2__EVAL_4;
  assign FormMicroOps__EVAL_108 = frontend__EVAL_96;
  assign ptw__EVAL_37 = core__EVAL_3;
  assign buffer_3__EVAL_30 = tlSlaveXbar__EVAL_9;
  assign coreXbar__EVAL_26 = filter__EVAL_42;
  assign rsource__EVAL_75 = _EVAL_75;
  assign dcache__EVAL_125 = ptw__EVAL_12;
  assign frontend__EVAL_63 = fragmenter__EVAL_27;
  assign tlMasterXbar__EVAL_52 = filter__EVAL_0;
  assign InstructionQueue__EVAL_86 = FormMicroOps__EVAL_103;
  assign ptw__EVAL_49 = core__EVAL_262;
  assign dcache__EVAL_122 = ptw__EVAL_104;
  assign frontend__EVAL_24 = fragmenter__EVAL_11;
  assign rsource__EVAL_101 = _EVAL_19;
  assign tlMasterXbar__EVAL_37 = filter__EVAL_63;
  assign dcache__EVAL_96 = dcacheArb__EVAL_7;
  assign core__EVAL_80 = InstructionQueue__EVAL_61;
  assign dcacheArb__EVAL_44 = dcache__EVAL_75;
  assign dcache__EVAL_52 = dcacheArb__EVAL_12;
  assign InstructionQueue__EVAL_58 = FormMicroOps__EVAL_63;
  assign frontend__EVAL_130 = ptw__EVAL_168;
  assign core__EVAL_236 = InstructionQueue__EVAL_144;
  assign core__EVAL_190 = dcacheArb__EVAL_20;
  assign core__EVAL_45 = InstructionQueue__EVAL_85;
  assign filter__EVAL_17 = coreXbar__EVAL_5;
  assign dcacheArb__EVAL_47 = core__EVAL_69;
  assign InstructionQueue__EVAL_167 = FormMicroOps__EVAL_35;
  assign ptw__EVAL_105 = core__EVAL_253;
  assign tlMasterXbar__EVAL_75 = buffer_2__EVAL;
  assign frontend__EVAL_131 = core__EVAL_225;
  assign frontend__EVAL_32 = fragmenter__EVAL_22;
  assign dcache__EVAL_5 = coreXbar__EVAL_69;
  assign InstructionQueue__EVAL_7 = FormMicroOps__EVAL_134;
  assign InstructionQueue__EVAL_101 = FormMicroOps__EVAL_82;
  assign coreXbar__EVAL_34 = widget_1__EVAL_32;
  assign fragmenter__EVAL_3 = _EVAL_32;
  assign InstructionQueue__EVAL_89 = FormMicroOps__EVAL_135;
  assign FormMicroOps__EVAL_110 = frontend__EVAL_84;
  assign frontend__EVAL_37 = ptw__EVAL_118;
  assign dlsXbar__EVAL_37 = widget_1__EVAL_3;
  assign dcache__EVAL_8 = dcacheArb__EVAL_19;
  assign frontend__EVAL_70 = ptw__EVAL_174;
  assign ptw__EVAL_70 = core__EVAL_140;
  assign core__EVAL_274 = InstructionQueue__EVAL_109;
  assign coreXbar__EVAL_0 = filter__EVAL_43;
  assign dcacheArb__EVAL_61 = core__EVAL_245;
  assign frontend__EVAL_81 = ptw__EVAL_74;
  assign buffer_2__EVAL_10 = rsource__EVAL_18;
  assign core__EVAL_92 = InstructionQueue__EVAL_0;
  assign core__EVAL_220 = InstructionQueue__EVAL_4;
  assign ptw__EVAL_132 = core__EVAL_14;
  assign core__EVAL_4 = intXbar__EVAL;
  assign InstructionQueue__EVAL_23 = FormMicroOps__EVAL_125;
  assign InstructionQueue__EVAL_50 = _EVAL_32 | core__EVAL_276;
  assign frontend__EVAL_78 = ptw__EVAL_136;
  assign rsource__EVAL_93 = _EVAL_86;
  assign ptw__EVAL_141 = core__EVAL_200;
  assign core__EVAL_170 = InstructionQueue__EVAL_2;
  assign fragmenter__EVAL_25 = widget__EVAL_19;
  assign core__EVAL_234 = dcacheArb__EVAL_62;
  assign rsource__EVAL_34 = _EVAL_91;
  assign frontend__EVAL_54 = core__EVAL_201;
  assign dcache__EVAL_4 = ptw__EVAL_1;
  assign InstructionQueue__EVAL_103 = FormMicroOps__EVAL_30;
  assign dcacheArb__EVAL_23 = core__EVAL_85;
  assign coreXbar__EVAL_38 = dcache__EVAL_92;
  assign _EVAL_13 = rsource__EVAL_59;
  assign core__EVAL_259 = dcacheArb__EVAL_74;
  assign dcacheArb__EVAL_90 = dcache__EVAL_128;
  assign InstructionQueue__EVAL_161 = FormMicroOps__EVAL_141;
  assign frontend__EVAL_113 = core__EVAL_276;
  assign widget__EVAL_21 = tlSlaveXbar__EVAL_35;
  assign core__EVAL_202 = InstructionQueue__EVAL_145;
  assign rsource__EVAL_22 = buffer_2__EVAL_41;
  assign frontend__EVAL_129 = core__EVAL_209;
  assign tlSlaveXbar__EVAL_28 = buffer_3__EVAL_37;
  assign core__EVAL_137 = InstructionQueue__EVAL_6;
  assign FormMicroOps__EVAL_91 = core__EVAL_128;
  assign widget__EVAL_26 = fragmenter__EVAL_19;
  assign coreXbar__EVAL_6 = dcache__EVAL_65;
  assign core__EVAL_31 = InstructionQueue__EVAL_162;
  assign buffer_2__EVAL_15 = rsource__EVAL_25;
  assign core__EVAL_169 = InstructionQueue__EVAL_118;
  assign rsource__EVAL_41 = _EVAL_61;
  assign ptw__EVAL_125 = core__EVAL_211;
  assign rsink__EVAL_8 = buffer_3__EVAL_33;
  assign rsink__EVAL_9 = _EVAL_98;
  assign buffer_2__EVAL_2 = tlMasterXbar__EVAL_65;
  assign buffer_2__EVAL_3 = rsource__EVAL_32;
  assign dcacheArb__EVAL_42 = dcache__EVAL_44;
  assign fragmenter_1__EVAL_14 = buffer_1__EVAL_4;
  assign buffer_1__EVAL_16 = dlsXbar__EVAL_34;
  assign _EVAL_52 = rsource__EVAL_51;
  assign rsink__EVAL_57 = buffer_3__EVAL_35;
  assign widget__EVAL_17 = tlSlaveXbar__EVAL_39;
  assign rsink__EVAL_14 = _EVAL_83;
  assign dcache__EVAL_58 = ptw__EVAL_24;
  assign dcache__EVAL_107 = coreXbar__EVAL_41;
  assign frontend__EVAL_90 = ptw__EVAL_63;
  assign dcacheArb__EVAL_29 = dcache__EVAL_105;
  assign FormMicroOps__EVAL_43 = frontend__EVAL_86;
  assign InstructionQueue__EVAL_71 = FormMicroOps__EVAL_114;
  assign core__EVAL_174 = dcacheArb__EVAL_27;
  assign dcache__EVAL_89 = ptw__EVAL_157;
  assign rsource__EVAL_44 = _EVAL_72;
  assign frontend__EVAL_48 = FormMicroOps__EVAL_34;
  assign _EVAL_33 = rsource__EVAL_46;
  assign ptw__EVAL_156 = core__EVAL_264;
  assign frontend__EVAL_74 = ptw__EVAL_82;
  assign widget__EVAL_13 = fragmenter__EVAL_26;
  assign core__EVAL_96 = InstructionQueue__EVAL_69;
  assign tlSlaveXbar__EVAL_45 = buffer_3__EVAL_26;
  assign intXbar__EVAL_5 = intsink_1__EVAL_3;
  assign frontend__EVAL_100 = ptw__EVAL_116;
  assign core__EVAL_57 = InstructionQueue__EVAL_81;
  assign core__EVAL_24 = dcacheArb__EVAL_10;
  assign fragmenter__EVAL_4 = frontend__EVAL_107;
  assign FormMicroOps__EVAL_136 = frontend__EVAL_61;
  assign intsink__EVAL_0 = _EVAL_100;
  assign InstructionQueue__EVAL_184 = FormMicroOps__EVAL_109;
  assign coreXbar__EVAL_82 = dcache__EVAL_126;
  assign InstructionQueue__EVAL_102 = FormMicroOps__EVAL_119;
  assign frontend__EVAL_83 = fragmenter__EVAL_13;
  assign dcache__EVAL_112 = coreXbar__EVAL_63;
  assign ptw__EVAL_28 = core__EVAL_189;
  assign dcacheArb__EVAL_45 = core__EVAL_248;
  assign dcacheArb__EVAL_56 = core__EVAL_167;
  assign frontend__EVAL_43 = buffer__EVAL_4;
  assign InstructionQueue__EVAL_147 = FormMicroOps__EVAL_70;
  assign frontend__EVAL_10 = buffer__EVAL_11;
  assign buffer_2__EVAL_48 = rsource__EVAL_55;
  assign frontend__EVAL_117 = ptw__EVAL_23;
  assign coreXbar__EVAL_79 = dcache__EVAL_103;
  assign core__EVAL_20 = InstructionQueue__EVAL_20;
  assign frontend__EVAL_13 = ptw__EVAL_94;
  assign buffer_2__EVAL_51 = tlMasterXbar__EVAL_27;
  assign buffer_2__EVAL_14 = tlMasterXbar__EVAL_43;
  assign rsource__EVAL_61 = _EVAL_64;
  assign ptw__EVAL_99 = core__EVAL_161;
  assign intsink_2__EVAL = _EVAL_100;
  assign dcache__EVAL_7 = ptw__EVAL_18;
  assign buffer_1__EVAL_7 = fragmenter_1__EVAL_10;
  assign core__EVAL_121 = InstructionQueue__EVAL_171;
  assign filter__EVAL_6 = coreXbar__EVAL_40;
  assign tlMasterXbar__EVAL_68 = buffer_2__EVAL_49;
  assign core__EVAL_32 = InstructionQueue__EVAL_155;
  assign filter__EVAL_12 = coreXbar__EVAL_62;
  assign dcache__EVAL_2 = ptw__EVAL_130;
  assign widget__EVAL_4 = tlSlaveXbar__EVAL_43;
  assign core__EVAL_64 = InstructionQueue__EVAL_125;
  assign rsink__EVAL_52 = _EVAL_36;
  assign _EVAL_95 = rsink__EVAL_38;
  assign buffer_3__EVAL_38 = rsink__EVAL_16;
  assign FormMicroOps__EVAL_12 = frontend__EVAL_125;
  assign coreXbar__EVAL_17 = dcache__EVAL_41;
  assign buffer__EVAL_7 = tlMasterXbar__EVAL_78;
  assign dcacheArb__EVAL_22 = dcache__EVAL_149;
  assign dcacheArb__EVAL_82 = dcache__EVAL_31;
  assign dcacheArb__EVAL_77 = dcache__EVAL_35;
  assign InstructionQueue__EVAL_80 = FormMicroOps__EVAL_62;
  assign core__EVAL_133 = dcacheArb__EVAL_17;
  assign coreXbar__EVAL_36 = filter__EVAL_7;
  assign InstructionQueue__EVAL_97 = FormMicroOps__EVAL_5;
  assign core__EVAL_277 = intXbar__EVAL_0;
  assign frontend__EVAL_109 = ptw__EVAL_134;
  assign filter__EVAL_66 = coreXbar__EVAL_78;
  assign frontend__EVAL_29 = ptw__EVAL_107;
  assign dcache__EVAL_90 = coreXbar__EVAL_14;
  assign core__EVAL_179 = InstructionQueue__EVAL_8;
  assign FormMicroOps__EVAL_31 = core__EVAL_231;
  assign InstructionQueue__EVAL_153 = FormMicroOps__EVAL_54;
  assign frontend__EVAL_121 = fragmenter__EVAL_28;
  assign dcache__EVAL_14 = coreXbar__EVAL_10;
  assign fragmenter_1__EVAL_22 = dls__EVAL_2;
  assign frontend__EVAL_64 = ptw__EVAL_86;
  assign coreXbar__EVAL_9 = widget_1__EVAL_18;
  assign tlMasterXbar__EVAL_22 = filter__EVAL_28;
  assign core__EVAL_22 = dcacheArb__EVAL_3;
  assign FormMicroOps__EVAL_6 = core__EVAL_82;
  assign ptw__EVAL_114 = core__EVAL_257;
  assign ptw__EVAL_73 = core__EVAL_113;
  assign rsource__EVAL_88 = _EVAL_7;
  assign FormMicroOps__EVAL_90 = core__EVAL_223;
  assign InstructionQueue__EVAL_117 = FormMicroOps__EVAL_158;
  assign core__EVAL_146 = dcacheArb__EVAL_50;
  assign _EVAL_105 = rsource__EVAL_16;
  assign dcache__EVAL_26 = ptw__EVAL_50;
  assign dcache__EVAL_81 = ptw__EVAL_66;
  assign dcache__EVAL_109 = ptw__EVAL_129;
  assign FormMicroOps__EVAL_92 = frontend__EVAL_75;
  assign ptw__EVAL_83 = core__EVAL_12;
  assign dcache__EVAL_40 = ptw__EVAL_61;
  assign tlMasterXbar__EVAL_13 = buffer_2__EVAL_20;
  assign frontend__EVAL_44 = _EVAL_32;
  assign ptw__EVAL_59 = core__EVAL_124;
  assign _EVAL_69 = rsource__EVAL_83;
  assign FormMicroOps__EVAL_48 = core__EVAL_30;
  assign _EVAL_92 = rsink__EVAL_33;
  assign FormMicroOps__EVAL_61 = frontend__EVAL_124;
  assign rsink__EVAL_51 = buffer_3__EVAL_19;
  assign dcache__EVAL_93 = ptw__EVAL_90;
  assign buffer_1__EVAL_26 = fragmenter_1__EVAL_24;
  assign rsource__EVAL_104 = buffer_2__EVAL_66;
  assign buffer_2__EVAL_58 = rsource__EVAL_90;
  assign rsink__EVAL_6 = buffer_3__EVAL_24;
  assign tlSlaveXbar__EVAL_49 = dlsXbar__EVAL_30;
  assign coreXbar__EVAL_33 = dcache__EVAL_80;
  assign dcache__EVAL_45 = ptw__EVAL_158;
  assign _EVAL_23 = rsink__EVAL_44;
  assign InstructionQueue__EVAL_41 = FormMicroOps__EVAL_80;
  assign ptw__EVAL_147 = core__EVAL_155;
  assign dcacheArb__EVAL_60 = dcache__EVAL_24;
  assign frontend__EVAL_6 = ptw__EVAL_40;
  assign InstructionQueue__EVAL_110 = FormMicroOps__EVAL_118;
  assign rsource__EVAL_11 = _EVAL_41;
  assign buffer_2__EVAL_19 = rsource__EVAL_87;
  assign _EVAL_43 = rsink__EVAL_37;
  assign FormMicroOps__EVAL_13 = frontend__EVAL_126;
  assign ptw__EVAL_178 = core__EVAL_103;
  assign filter__EVAL_4 = coreXbar__EVAL_59;
  assign fragmenter_1__EVAL_26 = buffer_1__EVAL_21;
  assign dlsXbar__EVAL_12 = tlSlaveXbar__EVAL_29;
  assign core__EVAL_163 = dcacheArb__EVAL_66;
  assign InstructionQueue__EVAL_62 = FormMicroOps__EVAL_123;
  assign buffer_2__EVAL_55 = tlMasterXbar__EVAL_39;
  assign widget_1__EVAL_12 = coreXbar__EVAL_87;
  assign ptw__EVAL_0 = core__EVAL_279;
  assign dcacheArb__EVAL_75 = dcache__EVAL_33;
  assign intsink_1__EVAL_0 = _EVAL_100;
  assign ptw__EVAL_2 = _EVAL_100;
  assign coreXbar__EVAL_73 = filter__EVAL_15;
  assign InstructionQueue__EVAL_48 = FormMicroOps__EVAL_41;
  assign InstructionQueue__EVAL_76 = FormMicroOps__EVAL_155;
  assign dcache__EVAL_38 = coreXbar__EVAL_43;
  assign rsink__EVAL_42 = _EVAL_59;
  assign InstructionQueue__EVAL_68 = FormMicroOps__EVAL_81;
  assign fragmenter_1__EVAL_6 = buffer_1__EVAL_27;
  assign tlMasterXbar__EVAL_82 = buffer__EVAL_3;
  assign _EVAL_71 = rsource__EVAL_9;
  assign InstructionQueue__EVAL_51 = FormMicroOps__EVAL_133;
  assign dlsXbar__EVAL_6 = widget_1__EVAL_30;
  assign ptw__EVAL_96 = core__EVAL_195;
  assign tlSlaveXbar__EVAL_2 = buffer_3__EVAL_6;
  assign buffer_2__EVAL_56 = tlMasterXbar__EVAL_2;
  assign core__EVAL_250 = InstructionQueue__EVAL_121;
  assign core__EVAL_29 = dcacheArb__EVAL_21;
  assign ptw__EVAL_5 = core__EVAL;
  assign ptw__EVAL_43 = core__EVAL_145;
  assign frontend__EVAL_85 = fragmenter__EVAL_6;
  assign InstructionQueue__EVAL_151 = FormMicroOps__EVAL_128;
  assign core__EVAL_78 = InstructionQueue__EVAL_34;
  assign rsource__EVAL_77 = _EVAL_42;
  assign dlsXbar__EVAL_3 = tlSlaveXbar__EVAL_30;
  assign dcache__EVAL_117 = dcacheArb__EVAL_28;
  assign buffer_2__EVAL_50 = tlMasterXbar__EVAL_58;
  assign buffer_2__EVAL_0 = tlMasterXbar__EVAL_25;
  assign _EVAL_40 = rsource__EVAL_97;
  assign frontend__EVAL_89 = core__EVAL_263;
  assign FormMicroOps__EVAL_27 = core__EVAL_273;
  assign rsource__EVAL_23 = buffer_2__EVAL_63;
  assign _EVAL_34 = rsource__EVAL_81;
  assign coreXbar__EVAL_35 = filter__EVAL_18;
  assign core__EVAL_255 = dcacheArb__EVAL_5;
  assign buffer_3__EVAL_15 = rsink__EVAL_19;
  assign FormMicroOps__EVAL_8 = frontend__EVAL_49;
  assign core__EVAL_237 = InstructionQueue__EVAL_182;
  assign core__EVAL_183 = InstructionQueue__EVAL_3;
  assign fragmenter_1__EVAL_15 = _EVAL_32;
  assign _EVAL_4 = rsource__EVAL_98;
  assign frontend__EVAL = _EVAL_38;
  assign ptw__EVAL_35 = core__EVAL_61;
  assign buffer_2__EVAL_61 = tlMasterXbar__EVAL_5;
  assign tlMasterXbar__EVAL_28 = filter__EVAL_16;
  assign FormMicroOps__EVAL_56 = core__EVAL_217;
  assign filter__EVAL_13 = coreXbar__EVAL_66;
  assign fragmenter_1__EVAL_25 = buffer_1__EVAL_31;
  assign InstructionQueue__EVAL_150 = FormMicroOps__EVAL_115;
  assign dcache__EVAL_87 = ptw__EVAL_45;
  assign rsource__EVAL_21 = _EVAL_107;
  assign dcache__EVAL_36 = coreXbar__EVAL_72;
  assign InstructionQueue__EVAL_32 = _EVAL_100;
  assign rsink__EVAL_40 = _EVAL_89;
  assign frontend__EVAL_39 = core__EVAL_41;
  assign filter__EVAL_8 = tlMasterXbar__EVAL_10;
  assign fragmenter__EVAL_23 = frontend__EVAL_110;
  assign frontend__EVAL_68 = ptw__EVAL_171;
  assign ptw__EVAL_101 = _EVAL_32;
  assign dls__EVAL_0 = fragmenter_1__EVAL_1;
  assign frontend__EVAL_30 = core__EVAL_192;
  assign core__EVAL_2 = InstructionQueue__EVAL_77;
  assign dcacheArb__EVAL_70 = dcache__EVAL_127;
  assign buffer_3__EVAL_23 = tlSlaveXbar__EVAL_8;
  assign dcacheArb__EVAL_11 = dcache__EVAL_119;
  assign core__EVAL_226 = InstructionQueue__EVAL_123;
  assign InstructionQueue__EVAL_137 = FormMicroOps__EVAL_71;
  assign dcacheArb__EVAL_41 = dcache__EVAL_84;
  assign FormMicroOps__EVAL_145 = core__EVAL_42;
  assign tlSlaveXbar__EVAL_15 = _EVAL_32;
  assign _EVAL = rsource__EVAL_95;
  assign frontend__EVAL_57 = _EVAL_100;
  assign InstructionQueue__EVAL_157 = FormMicroOps__EVAL_120;
  assign dcacheArb__EVAL_40 = core__EVAL_109;
  assign rsource__EVAL_35 = _EVAL_78;
  assign _EVAL_117 = rsink__EVAL_53;
  assign InstructionQueue__EVAL_44 = FormMicroOps__EVAL_149;
  assign tlSlaveXbar__EVAL_44 = dlsXbar__EVAL_22;
  assign tlSlaveXbar__EVAL_18 = dlsXbar__EVAL_0;
  assign dcacheArb__EVAL_0 = dcache__EVAL_146;
  assign InstructionQueue__EVAL_63 = FormMicroOps__EVAL_88;
  assign filter__EVAL_49 = _EVAL_32;
  assign ptw__EVAL_8 = core__EVAL_53;
  assign widget_1__EVAL_5 = coreXbar__EVAL_3;
  assign core__EVAL_261 = dcacheArb__EVAL;
  assign widget_1__EVAL_21 = dlsXbar__EVAL_41;
  assign filter__EVAL_60 = coreXbar__EVAL_45;
  assign coreXbar__EVAL_24 = _EVAL_32;
  assign dcacheArb__EVAL_18 = dcache__EVAL_143;
  assign buffer_1__EVAL_18 = dlsXbar__EVAL_10;
  assign buffer_3__EVAL_29 = rsink__EVAL_31;
  assign fragmenter__EVAL_10 = widget__EVAL_6;
  assign fragmenter_1__EVAL_7 = buffer_1__EVAL_13;
  assign core__EVAL_91 = InstructionQueue__EVAL_74;
  assign coreXbar__EVAL_68 = filter__EVAL_46;
  assign InstructionQueue__EVAL_87 = FormMicroOps__EVAL_22;
  assign dcache__EVAL_72 = _EVAL_100;
  assign frontend__EVAL_11 = core__EVAL_193;
  assign FormMicroOps__EVAL_29 = frontend__EVAL_25;
  assign fragmenter__EVAL_14 = frontend__EVAL_133;
  assign widget_1__EVAL_15 = coreXbar__EVAL_19;
  assign buffer_2__EVAL_72 = _EVAL_32;
  assign core__EVAL_213 = InstructionQueue__EVAL_84;
  assign FormMicroOps__EVAL_60 = core__EVAL_173;
  assign filter__EVAL_58 = coreXbar__EVAL_65;
  assign buffer_3__EVAL_9 = tlSlaveXbar__EVAL_41;
  assign FormMicroOps__EVAL_139 = core__EVAL_17;
  assign frontend__EVAL_82 = core__EVAL_18;
  assign frontend__EVAL_105 = ptw__EVAL_127;
  assign FormMicroOps__EVAL_47 = frontend__EVAL_106;
  assign fragmenter__EVAL_17 = _EVAL_100;
  assign frontend__EVAL_3 = ptw__EVAL_39;
  assign core__EVAL_242 = InstructionQueue__EVAL_40;
  assign rsink__EVAL_0 = _EVAL_22;
  assign coreXbar__EVAL_21 = filter__EVAL_20;
  assign dcache__EVAL_22 = ptw__EVAL_117;
  assign ptw__EVAL_109 = core__EVAL_160;
  assign tlMasterXbar__EVAL_29 = buffer_2__EVAL_5;
  assign coreXbar__EVAL_56 = dcache__EVAL_13;
  assign frontend__EVAL_51 = FormMicroOps__EVAL_46;
  assign rsink__EVAL_46 = _EVAL_12;
  assign core__EVAL_175 = dcacheArb__EVAL_15;
  assign rsource__EVAL_24 = _EVAL_111;
  assign dlsXbar__EVAL_40 = buffer_1__EVAL_32;
  assign dcache__EVAL_131 = ptw__EVAL_164;
  assign core__EVAL_115 = InstructionQueue__EVAL_93;
  assign tlMasterXbar__EVAL_67 = filter__EVAL_21;
  assign core__EVAL_216 = dcacheArb__EVAL_25;
  assign buffer_2__EVAL_32 = rsource__EVAL_45;
  assign widget__EVAL_20 = tlSlaveXbar__EVAL_12;
  assign FormMicroOps__EVAL_19 = core__EVAL_27;
  assign frontend__EVAL_15 = fragmenter__EVAL_21;
  assign InstructionQueue__EVAL_64 = FormMicroOps__EVAL_68;
  assign tlMasterXbar__EVAL_81 = buffer_2__EVAL_70;
  assign filter__EVAL_37 = coreXbar__EVAL_4;
  assign frontend__EVAL_112 = ptw__EVAL_111;
  assign frontend__EVAL_87 = ptw__EVAL_110;
  assign FormMicroOps__EVAL_107 = core__EVAL_239;
  assign coreXbar__EVAL_84 = dcache__EVAL_50;
  assign filter__EVAL_1 = tlMasterXbar__EVAL_45;
  assign tlSlaveXbar__EVAL_3 = widget__EVAL_22;
  assign core__EVAL_71 = InstructionQueue__EVAL_165;
  assign InstructionQueue__EVAL_16 = FormMicroOps__EVAL_3;
  assign dcache__EVAL_86 = coreXbar__EVAL_53;
  assign core__EVAL_63 = _EVAL_32;
  assign tlSlaveXbar__EVAL_27 = buffer_3__EVAL_7;
  assign buffer__EVAL_1 = tlMasterXbar__EVAL_36;
  assign FormMicroOps__EVAL_156 = core__EVAL_120;
  assign frontend__EVAL_71 = ptw__EVAL_124;
  assign tlMasterXbar__EVAL_4 = buffer_2__EVAL_65;
  assign dcacheArb__EVAL_80 = dcache__EVAL_129;
  assign coreXbar__EVAL_16 = dcache__EVAL_15;
  assign tlSlaveXbar__EVAL_20 = widget__EVAL_18;
  assign dlsXbar__EVAL_28 = tlSlaveXbar__EVAL_36;
  assign dcache__EVAL_69 = ptw__EVAL_22;
  assign FormMicroOps__EVAL_66 = _EVAL_32 | core__EVAL_276;
  assign rsource__EVAL_42 = _EVAL_32;
  assign InstructionQueue__EVAL_107 = FormMicroOps__EVAL_94;
  assign _EVAL_35 = rsource__EVAL_39;
  assign frontend__EVAL_114 = ptw__EVAL_14;
  assign frontend__EVAL_104 = ptw__EVAL_172;
  assign FormMicroOps__EVAL_9 = core__EVAL_7;
  assign dcache__EVAL_101 = ptw__EVAL_146;
  assign filter__EVAL_56 = tlMasterXbar__EVAL;
  assign fragmenter__EVAL = widget__EVAL_2;
  assign frontend__EVAL_9 = ptw__EVAL_68;
  assign dcache__EVAL_145 = coreXbar__EVAL_86;
  assign _EVAL_16 = rsource__EVAL_31;
  assign _EVAL_73 = rsource__EVAL_103;
  assign buffer_2__EVAL_7 = rsource__EVAL_91;
  assign frontend__EVAL_55 = ptw__EVAL_108;
  assign ptw__EVAL_121 = core__EVAL_52;
  assign widget_1__EVAL_25 = coreXbar__EVAL_81;
  assign ptw__EVAL_81 = core__EVAL_271;
  assign core__EVAL_87 = dcacheArb__EVAL_26;
  assign FormMicroOps__EVAL_142 = core__EVAL_100;
  assign dcache__EVAL_85 = ptw__EVAL_31;
  assign dcache__EVAL_9 = ptw__EVAL_100;
  assign dcache__EVAL_115 = ptw__EVAL_170;
  assign tlMasterXbar__EVAL_49 = buffer_2__EVAL_64;
  assign buffer_3__EVAL_10 = tlSlaveXbar__EVAL_33;
  assign rsource__EVAL_29 = buffer_2__EVAL_52;
  assign frontend__EVAL_19 = core__EVAL_65;
  assign core__EVAL_95 = frontend__EVAL_17;
  assign _EVAL_116 = rsource__EVAL_30;
  assign dcache__EVAL_135 = dcacheArb__EVAL_71;
  assign coreXbar__EVAL_29 = dcache__EVAL_57;
  assign ptw__EVAL_34 = core__EVAL_197;
  assign FormMicroOps__EVAL_152 = frontend__EVAL_102;
  assign dcache__EVAL_120 = ptw__EVAL_11;
  assign core__EVAL_212 = InstructionQueue__EVAL_53;
  assign _EVAL_118 = rsink__EVAL_7;
  assign coreXbar__EVAL_27 = dcache__EVAL_147;
  assign widget_1__EVAL_4 = dlsXbar__EVAL_33;
  assign widget__EVAL_23 = fragmenter__EVAL_0;
  assign core__EVAL_148 = InstructionQueue__EVAL_112;
  assign core__EVAL_84 = InstructionQueue__EVAL_183;
  assign InstructionQueue__EVAL_119 = FormMicroOps__EVAL_74;
  assign tlMasterXbar__EVAL_17 = filter__EVAL_5;
  assign buffer_3__EVAL_36 = rsink__EVAL_5;
  assign frontend__EVAL_92 = ptw__EVAL_6;
  assign buffer__EVAL_19 = _EVAL_100;
  assign rsink__EVAL_56 = buffer_3__EVAL_11;
  assign widget__EVAL_9 = _EVAL_100;
  assign InstructionQueue__EVAL_127 = FormMicroOps__EVAL_130;
  assign core__EVAL_164 = InstructionQueue__EVAL_66;
  assign buffer_3__EVAL_16 = rsink__EVAL_45;
  assign ptw__EVAL_67 = core__EVAL_136;
  assign frontend__EVAL_50 = ptw__EVAL_62;
  assign dls__EVAL_5 = fragmenter_1__EVAL_17;
  assign _EVAL_82 = rsource__EVAL_79;
  assign InstructionQueue__EVAL_10 = FormMicroOps__EVAL_37;
  assign core__EVAL_147 = dcacheArb__EVAL_59;
  assign filter__EVAL = coreXbar__EVAL_80;
  assign frontend__EVAL_4 = ptw__EVAL_19;
  assign core__EVAL_247 = InstructionQueue__EVAL_166;
  assign dcache__EVAL_114 = ptw__EVAL_53;
  assign intsink_1__EVAL_2 = _EVAL_9;
  assign _EVAL_114 = rsink__EVAL_24;
  assign buffer_1__EVAL_10 = fragmenter_1__EVAL_4;
  assign buffer__EVAL_10 = _EVAL_32;
  assign filter__EVAL_2 = coreXbar__EVAL_12;
  assign InstructionQueue__EVAL_168 = FormMicroOps__EVAL_116;
  assign InstructionQueue__EVAL_33 = FormMicroOps__EVAL_21;
  assign InstructionQueue__EVAL_156 = FormMicroOps__EVAL_97;
  assign core__EVAL_68 = InstructionQueue__EVAL_13;
  assign InstructionQueue__EVAL_100 = FormMicroOps__EVAL;
  assign _EVAL_108 = rsource__EVAL_65;
  assign coreXbar__EVAL_50 = filter__EVAL_26;
  assign dcache__EVAL_142 = ptw__EVAL_140;
  assign fragmenter__EVAL_24 = widget__EVAL_0;
  assign FormMicroOps__EVAL_100 = frontend__EVAL_31;
  assign InstructionQueue__EVAL_104 = FormMicroOps__EVAL_14;
  assign tlSlaveXbar__EVAL_26 = _EVAL_100;
  assign dcache__EVAL_124 = dcacheArb__EVAL_48;
  assign tlMasterXbar__EVAL_83 = _EVAL_32;
  assign dlsXbar__EVAL_17 = _EVAL_100;
  assign InstructionQueue__EVAL_14 = FormMicroOps__EVAL_4;
  assign tlMasterXbar__EVAL_70 = buffer_2__EVAL_59;
  assign tlSlaveXbar__EVAL_5 = dlsXbar__EVAL_38;
  assign filter__EVAL_64 = coreXbar__EVAL_64;
  assign frontend__EVAL_0 = ptw__EVAL_155;
  assign rsink__EVAL_12 = _EVAL_6;
  assign buffer_1__EVAL_29 = fragmenter_1__EVAL_12;
  assign InstructionQueue__EVAL_154 = FormMicroOps__EVAL_0;
  assign rsource__EVAL_70 = _EVAL_51;
  assign buffer_3__EVAL_18 = rsink__EVAL_28;
  assign frontend__EVAL_67 = ptw__EVAL_153;
  assign buffer_2__EVAL_30 = rsource__EVAL_38;
  assign rsource__EVAL_82 = buffer_2__EVAL_31;
  assign InstructionQueue__EVAL_116 = FormMicroOps__EVAL_106;
  assign ptw__EVAL_20 = core__EVAL_235;
  assign rsink__EVAL_27 = _EVAL_100;
  assign dcache__EVAL_137 = coreXbar__EVAL_75;
  assign coreXbar__EVAL_42 = widget_1__EVAL_10;
  assign InstructionQueue__EVAL_29 = FormMicroOps__EVAL_2;
  assign dcacheArb__EVAL_57 = core__EVAL_34;
  assign core__EVAL_184 = InstructionQueue__EVAL_22;
  assign frontend__EVAL_35 = ptw__EVAL_126;
  assign FormMicroOps__EVAL_147 = core__EVAL_243;
  assign buffer__EVAL_17 = frontend__EVAL_108;
  assign rsink__EVAL_49 = _EVAL_55;
  assign core__EVAL_141 = InstructionQueue__EVAL_79;
  assign fragmenter__EVAL_5 = widget__EVAL_14;
  assign dcache__EVAL_79 = ptw__EVAL_26;
  assign widget_1__EVAL_23 = coreXbar__EVAL_76;
  assign core__EVAL_25 = dcacheArb__EVAL_83;
  assign InstructionQueue__EVAL_169 = FormMicroOps__EVAL_38;
  assign buffer_2__EVAL_9 = tlMasterXbar__EVAL_66;
  assign frontend__EVAL_2 = core__EVAL_185;
  assign ptw__EVAL_21 = core__EVAL_240;
  assign fragmenter_1__EVAL_31 = buffer_1__EVAL_6;
  assign FormMicroOps__EVAL_144 = core__EVAL_19;
  assign InstructionQueue__EVAL_142 = FormMicroOps__EVAL_86;
  assign dcache__EVAL_132 = ptw__EVAL_151;
  assign _EVAL_97 = rsink__EVAL_54;
  assign fragmenter__EVAL_18 = frontend__EVAL_69;
  assign tlMasterXbar__EVAL_59 = buffer_2__EVAL_27;
  assign buffer_1__EVAL_9 = dlsXbar__EVAL_48;
  assign widget_1__EVAL_17 = _EVAL_32;
  assign FormMicroOps__EVAL_95 = frontend__EVAL_99;
  assign buffer_1__EVAL_0 = dlsXbar__EVAL_21;
  assign rsource__EVAL_74 = buffer_2__EVAL_34;
  assign dcache__EVAL_78 = ptw__EVAL_76;
  assign FormMicroOps__EVAL_117 = frontend__EVAL_62;
  assign FormMicroOps__EVAL_49 = core__EVAL_74;
  assign core__EVAL_191 = InstructionQueue__EVAL_9;
  assign ptw__EVAL = core__EVAL_46;
  assign buffer_2__EVAL_68 = tlMasterXbar__EVAL_63;
  assign InstructionQueue__EVAL_148 = FormMicroOps__EVAL_150;
  assign core__EVAL_104 = InstructionQueue__EVAL_124;
  assign ptw__EVAL_133 = core__EVAL_9;
  assign rsource__EVAL_33 = _EVAL_50;
  assign dls__EVAL_8 = fragmenter_1__EVAL;
  assign FormMicroOps__EVAL_25 = core__EVAL_221;
  assign rsource__EVAL_71 = buffer_2__EVAL_45;
  assign rsource__EVAL_56 = buffer_2__EVAL_36;
  assign InstructionQueue__EVAL_172 = FormMicroOps__EVAL_151;
  assign buffer_3__EVAL_27 = rsink__EVAL_20;
  assign tlSlaveXbar__EVAL_10 = buffer_3__EVAL_8;
  assign dcache__EVAL_139 = dcacheArb__EVAL_2;
  assign coreXbar__EVAL_11 = dcache__EVAL_134;
  assign FormMicroOps__EVAL_75 = frontend__EVAL_56;
  assign dlsXbar__EVAL_13 = widget_1__EVAL_2;
  assign rsource__EVAL_12 = buffer_2__EVAL_26;
  assign dcacheArb__EVAL_38 = core__EVAL_94;
  assign dcacheArb__EVAL_64 = dcache__EVAL;
  assign dls__EVAL_15 = fragmenter_1__EVAL_32;
  assign buffer_2__EVAL_53 = rsource__EVAL_94;
  assign coreXbar__EVAL_58 = filter__EVAL_27;
  assign filter__EVAL_45 = tlMasterXbar__EVAL_34;
  assign dcache__EVAL_27 = ptw__EVAL_167;
  assign tlSlaveXbar__EVAL = dlsXbar__EVAL_2;
  assign core__EVAL_156 = frontend__EVAL_22;
  assign _EVAL_113 = rsink__EVAL_2;
  assign frontend__EVAL_28 = ptw__EVAL_29;
  assign tlMasterXbar__EVAL_50 = filter__EVAL_3;
  assign dcacheArb__EVAL_52 = dcache__EVAL_48;
  assign core__EVAL_222 = InstructionQueue__EVAL_163;
  assign widget_1__EVAL_8 = coreXbar__EVAL_39;
  assign buffer__EVAL_2 = tlMasterXbar__EVAL_42;
  assign coreXbar__EVAL_7 = _EVAL_100;
  assign tlMasterXbar__EVAL_20 = filter__EVAL_36;
  assign dcache__EVAL_23 = ptw__EVAL_166;
  assign dcache__EVAL_18 = _EVAL_32;
  assign dls__EVAL_9 = fragmenter_1__EVAL_21;
  assign dcache__EVAL_118 = ptw__EVAL_138;
  assign InstructionQueue__EVAL_174 = FormMicroOps__EVAL_105;
  assign core__EVAL_108 = InstructionQueue__EVAL_57;
  assign core__EVAL_106 = InstructionQueue__EVAL_49;
  assign core__EVAL_265 = InstructionQueue__EVAL_45;
  assign dcacheArb__EVAL_34 = dcache__EVAL_32;
  assign _EVAL_17 = rsource__EVAL_1;
  assign buffer_1__EVAL_1 = _EVAL_100;
  assign core__EVAL_1 = InstructionQueue__EVAL_73;
  assign buffer_2__EVAL_54 = tlMasterXbar__EVAL_64;
  assign core__EVAL_171 = InstructionQueue__EVAL_91;
  assign dlsXbar__EVAL_32 = widget_1__EVAL_11;
  assign dcache__EVAL_0 = ptw__EVAL_139;
  assign frontend__EVAL_141 = core__EVAL_182;
  assign ptw__EVAL_64 = core__EVAL_86;
  assign InstructionQueue__EVAL_131 = FormMicroOps__EVAL_18;
  assign InstructionQueue__EVAL_164 = FormMicroOps__EVAL_50;
  assign buffer__EVAL_9 = tlMasterXbar__EVAL_55;
  assign intXbar__EVAL_4 = intsink__EVAL;
  assign dcache__EVAL_140 = ptw__EVAL_88;
  assign ptw__EVAL_56 = core__EVAL_135;
  assign rsink__EVAL_1 = _EVAL_39;
  assign frontend__EVAL_23 = ptw__EVAL_87;
  assign fragmenter_1__EVAL_19 = dls__EVAL_14;
  assign ptw__EVAL_162 = core__EVAL_112;
  assign tlMasterXbar__EVAL_44 = filter__EVAL_59;
  assign dcache__EVAL_74 = ptw__EVAL_30;
  assign InstructionQueue__EVAL_178 = FormMicroOps__EVAL_112;
  assign rsource__EVAL_7 = _EVAL_100;
  assign dls__EVAL_10 = fragmenter_1__EVAL_23;
  assign filter__EVAL_57 = tlMasterXbar__EVAL_62;
  assign rsink__EVAL_58 = _EVAL_101;
  assign InstructionQueue__EVAL_181 = FormMicroOps__EVAL_83;
  assign ptw__EVAL_142 = core__EVAL_149;
  assign buffer_2__EVAL_71 = tlMasterXbar__EVAL_16;
  assign ptw__EVAL_58 = core__EVAL_228;
  assign core__EVAL_36 = frontend__EVAL_72;
  assign buffer_3__EVAL_22 = rsink__EVAL_18;
  assign dcache__EVAL_99 = coreXbar__EVAL_85;
  assign filter__EVAL_69 = coreXbar__EVAL_71;
  assign _EVAL_103 = rsource__EVAL_14;
  assign dcache__EVAL_88 = ptw__EVAL_57;
  assign FormMicroOps__EVAL_127 = frontend__EVAL_79;
  assign buffer_3__EVAL_5 = tlSlaveXbar__EVAL_6;
  assign tlSlaveXbar__EVAL_25 = buffer_3__EVAL_31;
  assign dcache__EVAL_53 = ptw__EVAL_79;
  assign core__EVAL_134 = intXbar__EVAL_2;
  assign InstructionQueue__EVAL_115 = FormMicroOps__EVAL_7;
  assign filter__EVAL_32 = tlMasterXbar__EVAL_35;
  assign coreXbar__EVAL_18 = dcache__EVAL_46;
  assign ptw__EVAL_4 = core__EVAL_139;
  assign coreXbar__EVAL_22 = dcache__EVAL_123;
  assign InstructionQueue__EVAL_75 = FormMicroOps__EVAL_28;
  assign _EVAL_106 = rsource__EVAL;
  assign dcacheArb__EVAL_69 = dcache__EVAL_68;
  assign widget__EVAL_1 = fragmenter__EVAL_9;
  assign tlMasterXbar__EVAL_47 = buffer_2__EVAL_46;
  assign InstructionQueue__EVAL_114 = FormMicroOps__EVAL_20;
  assign dcache__EVAL_97 = ptw__EVAL_123;
  assign filter__EVAL_52 = coreXbar__EVAL_25;
  assign filter__EVAL_70 = tlMasterXbar__EVAL_11;
  assign _EVAL_85 = rsink__EVAL_55;
  assign InstructionQueue__EVAL_25 = FormMicroOps__EVAL_153;
  assign frontend__EVAL_101 = ptw__EVAL_41;
  assign core__EVAL_111 = dcacheArb__EVAL_76;
  assign _EVAL_49 = rsink__EVAL_25;
  assign _EVAL_110 = rsink__EVAL_36;
  assign dcache__EVAL_25 = ptw__EVAL_44;
  assign buffer_2__EVAL_11 = tlMasterXbar__EVAL_15;
  assign dcache__EVAL_106 = ptw__EVAL_137;
  assign buffer_3__EVAL_20 = tlSlaveXbar__EVAL_1;
  assign rsink__EVAL_29 = _EVAL_84;
  assign widget__EVAL_5 = tlSlaveXbar__EVAL_7;
  assign dcacheArb__EVAL_8 = dcache__EVAL_61;
  assign core__EVAL_76 = InstructionQueue__EVAL_52;
  assign rsink__EVAL_50 = _EVAL_53;
  assign frontend__EVAL_7 = ptw__EVAL_42;
  assign filter__EVAL_41 = tlMasterXbar__EVAL_38;
  assign buffer__EVAL_16 = tlMasterXbar__EVAL_41;
  assign rsource__EVAL_89 = buffer_2__EVAL_17;
  assign core__EVAL_105 = intXbar__EVAL_3;
  assign coreXbar__EVAL_28 = dcache__EVAL_76;
  assign InstructionQueue__EVAL_12 = FormMicroOps__EVAL_45;
  assign dcacheArb__EVAL_43 = dcache__EVAL_82;
  assign _EVAL_76 = rsource__EVAL_28;
  assign frontend__EVAL_58 = ptw__EVAL_97;
  assign filter__EVAL_9 = tlMasterXbar__EVAL_40;
  assign FormMicroOps__EVAL_26 = InstructionQueue__EVAL_176;
  assign frontend__EVAL_5 = ptw__EVAL_60;
  assign ptw__EVAL_33 = core__EVAL_83;
  assign widget__EVAL_16 = tlSlaveXbar__EVAL_17;
  assign buffer__EVAL_6 = tlMasterXbar__EVAL_30;
  assign InstructionQueue__EVAL_177 = FormMicroOps__EVAL_157;
  assign frontend__EVAL_38 = core__EVAL_43;
  assign tlMasterXbar__EVAL_71 = buffer_2__EVAL_12;
  assign dlsXbar__EVAL = buffer_1__EVAL_11;
  assign buffer_2__EVAL_25 = tlMasterXbar__EVAL_31;
  assign dcacheArb__EVAL_63 = core__EVAL_116;
  assign frontend__EVAL_16 = core__EVAL_33;
  assign tlMasterXbar__EVAL_76 = buffer_2__EVAL_28;
  assign tlSlaveXbar__EVAL_32 = dlsXbar__EVAL_46;
  assign frontend__EVAL_33 = ptw__EVAL_54;
  assign core__EVAL_186 = InstructionQueue__EVAL_138;
  assign core__EVAL_73 = InstructionQueue__EVAL_129;
  assign dls__EVAL_4 = fragmenter_1__EVAL_29;
  assign InstructionQueue__EVAL_31 = FormMicroOps__EVAL_111;
  assign core__EVAL_158 = InstructionQueue__EVAL_128;
  assign rsource__EVAL_60 = buffer_2__EVAL_43;
  assign frontend__EVAL_60 = ptw__EVAL_3;
  assign _EVAL_56 = rsink__EVAL_48;
  assign InstructionQueue__EVAL_5 = FormMicroOps__EVAL_84;
  assign _EVAL_25 = rsource__EVAL_40;
  assign core__EVAL_39 = InstructionQueue__EVAL_140;
  assign ptw__EVAL_148 = core__EVAL_143;
  assign coreXbar__EVAL_23 = dcache__EVAL_6;
  assign ptw__EVAL_161 = core__EVAL_132;
  assign rsource__EVAL_3 = buffer_2__EVAL_6;
  assign rsink__EVAL_32 = buffer_3__EVAL_4;
  assign fragmenter_1__EVAL_13 = dls__EVAL_16;
  assign fragmenter_1__EVAL_16 = dls__EVAL_3;
  assign filter__EVAL_39 = _EVAL_100;
  assign widget__EVAL_3 = fragmenter__EVAL_2;
  assign frontend__EVAL_59 = ptw__EVAL_36;
  assign rsource__EVAL_17 = buffer_2__EVAL_47;
  assign frontend__EVAL_45 = core__EVAL_177;
  assign buffer__EVAL_12 = frontend__EVAL_66;
  assign InstructionQueue__EVAL_175 = FormMicroOps__EVAL_69;
  assign frontend__EVAL_52 = ptw__EVAL_135;
  assign FormMicroOps__EVAL_72 = core__EVAL_8;
  assign dlsXbar__EVAL_43 = tlSlaveXbar__EVAL_38;
  assign rsink__EVAL_60 = buffer_3__EVAL_34;
  assign buffer_1__EVAL_2 = dlsXbar__EVAL_27;
  assign InstructionQueue__EVAL_19 = core__EVAL_254;
  assign rsource__EVAL_106 = buffer_2__EVAL_62;
  assign _EVAL_62 = rsource__EVAL_5;
  assign dcacheArb__EVAL_1 = dcache__EVAL_34;
  assign core__EVAL_180 = InstructionQueue__EVAL_133;
  assign intXbar__EVAL_1 = intsink_1__EVAL;
  assign InstructionQueue__EVAL_54 = FormMicroOps__EVAL_101;
  assign tlMasterXbar__EVAL_79 = filter__EVAL_47;
  assign rsource__EVAL_100 = buffer_2__EVAL_23;
  assign rsource__EVAL_68 = _EVAL_26;
  assign dcache__EVAL_21 = ptw__EVAL_93;
  assign core__EVAL_6 = InstructionQueue__EVAL_141;
  assign core__EVAL_272 = InstructionQueue__EVAL_111;
  assign rsource__EVAL_105 = _EVAL_112;
  assign tlMasterXbar__EVAL_80 = _EVAL_100;
  assign dcacheArb__EVAL_46 = dcache__EVAL_42;
  assign widget_1__EVAL_1 = dlsXbar__EVAL_18;
  assign frontend__EVAL_139 = core__EVAL_151;
  assign dcache__EVAL_56 = dcacheArb__EVAL_85;
  assign FormMicroOps__EVAL_102 = core__EVAL_187;
  assign dlsXbar__EVAL_1 = widget_1__EVAL_20;
  assign ptw__EVAL_27 = core__EVAL_194;
  assign InstructionQueue__EVAL_55 = FormMicroOps__EVAL_129;
  assign InstructionQueue__EVAL_158 = FormMicroOps__EVAL_85;
  assign _EVAL_87 = rsource__EVAL_47;
  assign _EVAL_58 = rsink__EVAL_23;
  assign frontend__EVAL_12 = core__EVAL_99;
  assign _EVAL_60 = rsink__EVAL_34;
  assign frontend__EVAL_27 = ptw__EVAL_150;
  assign dcache__EVAL_66 = coreXbar__EVAL_74;
  assign buffer_2__EVAL_42 = rsource__EVAL_76;
  assign InstructionQueue__EVAL_37 = FormMicroOps__EVAL_17;
  assign FormMicroOps__EVAL_122 = frontend__EVAL_26;
  assign dcacheArb__EVAL_49 = core__EVAL_118;
  assign tlSlaveXbar__EVAL_16 = buffer_3__EVAL_3;
  assign coreXbar__EVAL_77 = filter__EVAL_54;
  assign dcacheArb__EVAL_36 = core__EVAL_62;
  assign InstructionQueue__EVAL_130 = FormMicroOps__EVAL_36;
  assign dcache__EVAL_12 = ptw__EVAL_120;
  assign dcache__EVAL_63 = ptw__EVAL_92;
  assign fragmenter__EVAL_16 = widget__EVAL_15;
  assign InstructionQueue__EVAL_47 = FormMicroOps__EVAL_137;
  assign widget_1__EVAL_13 = dlsXbar__EVAL_11;
  assign InstructionQueue__EVAL_126 = FormMicroOps__EVAL_146;
  assign frontend__EVAL_142 = core__EVAL_117;
  assign core__EVAL_214 = InstructionQueue__EVAL_90;
  assign intXbar__EVAL_6 = intsink_2__EVAL_1;
  assign ptw__EVAL_144 = core__EVAL_131;
  assign core__EVAL_270 = _EVAL_38;
  assign intsink_1__EVAL_1 = _EVAL_47;
  assign dcache__EVAL_98 = ptw__EVAL_75;
  assign filter__EVAL_22 = coreXbar__EVAL_15;
  assign rsource__EVAL_15 = _EVAL_45;
  assign InstructionQueue__EVAL = FormMicroOps__EVAL_124;
  assign core__EVAL_153 = InstructionQueue__EVAL_18;
  assign frontend__EVAL_132 = buffer__EVAL_18;
  assign rsource__EVAL_13 = _EVAL_74;
  assign dls__EVAL_1 = _EVAL_100;
  assign InstructionQueue__EVAL_88 = FormMicroOps__EVAL_96;
  assign _EVAL_44 = rsink__EVAL;
  assign ptw__EVAL_69 = core__EVAL_199;
  assign core__EVAL_58 = InstructionQueue__EVAL_96;
  assign frontend__EVAL_8 = ptw__EVAL_80;
  assign core__EVAL_260 = InstructionQueue__EVAL_179;
  assign coreXbar__EVAL_88 = filter__EVAL_67;
  assign frontend__EVAL_42 = ptw__EVAL_175;
  assign _EVAL_5 = rsink__EVAL_3;
  assign InstructionQueue__EVAL_28 = FormMicroOps__EVAL_23;
  assign tlMasterXbar__EVAL_51 = buffer_2__EVAL_24;
  assign dls__EVAL_11 = fragmenter_1__EVAL_11;
  assign InstructionQueue__EVAL_60 = core__EVAL_129;
  assign tlMasterXbar__EVAL_77 = filter__EVAL_68;
  assign FormMicroOps__EVAL_33 = frontend__EVAL_53;
  assign buffer_2__EVAL_21 = tlMasterXbar__EVAL_1;
  assign tlMasterXbar__EVAL_26 = buffer_2__EVAL_29;
  assign fragmenter__EVAL_1 = widget__EVAL_27;
  assign dcache__EVAL_51 = ptw__EVAL_65;
  assign frontend__EVAL_137 = fragmenter__EVAL_20;
  assign tlSlaveXbar__EVAL_0 = buffer_3__EVAL_25;
  assign _EVAL_81 = rsource__EVAL_99;
  assign FormMicroOps__EVAL_57 = core__EVAL_207;
  assign InstructionQueue__EVAL_11 = FormMicroOps__EVAL_40;
  assign dlsXbar__EVAL_4 = tlSlaveXbar__EVAL_4;
  assign buffer_3__EVAL_17 = rsink__EVAL_11;
  assign InstructionQueue__EVAL_72 = FormMicroOps__EVAL_59;
  assign FormMicroOps__EVAL_79 = core__EVAL_26;
  assign coreXbar__EVAL_13 = widget_1__EVAL_0;
  assign core__EVAL_98 = InstructionQueue__EVAL_78;
  assign InstructionQueue__EVAL_82 = FormMicroOps__EVAL_131;
  assign core__EVAL_47 = dcacheArb__EVAL_16;
  assign core__EVAL_233 = dcacheArb__EVAL_73;
  assign filter__EVAL_48 = coreXbar__EVAL_47;
  assign dcache__EVAL_55 = ptw__EVAL_145;
  assign ptw__EVAL_112 = core__EVAL_66;
  assign InstructionQueue__EVAL_36 = FormMicroOps__EVAL_55;
  assign frontend__EVAL_65 = core__EVAL_56;
  assign FormMicroOps__EVAL_77 = core__EVAL_0;
  assign buffer_3__EVAL_21 = rsink__EVAL_26;
  assign frontend__EVAL_73 = ptw__EVAL_152;
  assign InstructionQueue__EVAL_1 = FormMicroOps__EVAL_15;
  assign dlsXbar__EVAL_45 = widget_1__EVAL;
  assign widget_1__EVAL_6 = dlsXbar__EVAL_9;
  assign InstructionQueue__EVAL_95 = FormMicroOps__EVAL_65;
  assign core__EVAL_204 = InstructionQueue__EVAL_113;
  assign rsource__EVAL_50 = _EVAL_54;
  assign InstructionQueue__EVAL_108 = FormMicroOps__EVAL_76;
  assign rsink__EVAL_59 = buffer_3__EVAL;
  assign dcacheArb__EVAL_4 = dcache__EVAL_136;
  assign tlMasterXbar__EVAL_56 = filter__EVAL_40;
  assign dcache__EVAL_20 = coreXbar__EVAL_32;
  assign dcache__EVAL_113 = ptw__EVAL_48;
  assign dcacheArb__EVAL_24 = dcache__EVAL_110;
  assign _EVAL_109 = rsource__EVAL_73;
  assign core__EVAL_205 = InstructionQueue__EVAL_160;
  assign tlMasterXbar__EVAL_23 = filter__EVAL_55;
  assign dcache__EVAL_144 = ptw__EVAL_149;
  assign buffer_3__EVAL_32 = tlSlaveXbar__EVAL_14;
  assign FormMicroOps__EVAL_32 = core__EVAL_252;
  assign widget_1__EVAL_7 = coreXbar__EVAL_52;
  assign buffer_2__EVAL_67 = tlMasterXbar__EVAL_18;
  assign frontend__EVAL_118 = core__EVAL_275;
  assign buffer_2__EVAL_38 = rsource__EVAL_53;
  assign buffer_1__EVAL_3 = dlsXbar__EVAL_25;
  assign rsink__EVAL_10 = _EVAL_70;
  assign widget__EVAL_25 = fragmenter__EVAL_15;
  assign dls__EVAL = _EVAL_32;
  assign fragmenter__EVAL_8 = frontend__EVAL_76;
  assign _EVAL_20 = rsource__EVAL_43;
  assign widget_1__EVAL_26 = _EVAL_100;
  assign tlSlaveXbar__EVAL_48 = widget__EVAL_8;
  assign rsource__EVAL_66 = _EVAL_21;
  assign dcache__EVAL_116 = ptw__EVAL_15;
endmodule
