//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_29(
  output        _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  output [10:0] _EVAL_2,
  output [3:0]  _EVAL_3,
  input  [10:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  output [3:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  output [3:0]  _EVAL_9,
  input         _EVAL_10,
  output        _EVAL_11,
  input  [7:0]  _EVAL_12,
  output        _EVAL_13,
  input  [10:0] _EVAL_14,
  input  [3:0]  _EVAL_15,
  output [10:0] _EVAL_16,
  input  [10:0] _EVAL_17,
  output [1:0]  _EVAL_18,
  input         _EVAL_19,
  output [3:0]  _EVAL_20,
  input  [3:0]  _EVAL_21,
  input         _EVAL_22,
  input  [2:0]  _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output [31:0] _EVAL_26,
  input  [7:0]  _EVAL_27,
  input         _EVAL_28,
  output [2:0]  _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  output [1:0]  _EVAL_32,
  output [3:0]  _EVAL_33,
  input  [2:0]  _EVAL_34,
  input         _EVAL_35,
  input  [3:0]  _EVAL_36,
  input  [31:0] _EVAL_37,
  output [30:0] _EVAL_38,
  output        _EVAL_39,
  input  [30:0] _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  output [3:0]  _EVAL_43,
  input  [10:0] _EVAL_44,
  output [2:0]  _EVAL_45,
  input  [3:0]  _EVAL_46,
  input  [3:0]  _EVAL_47,
  output        _EVAL_48,
  output [1:0]  _EVAL_49,
  input  [1:0]  _EVAL_50,
  input  [2:0]  _EVAL_51,
  output [7:0]  _EVAL_52,
  output [2:0]  _EVAL_53,
  output [1:0]  _EVAL_54,
  output [30:0] _EVAL_55,
  input  [1:0]  _EVAL_56,
  output [2:0]  _EVAL_57,
  input  [1:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  input         _EVAL_60,
  output [10:0] _EVAL_61,
  input  [2:0]  _EVAL_62,
  input  [3:0]  _EVAL_63,
  input  [30:0] _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  output [2:0]  _EVAL_67,
  input         _EVAL_68,
  input  [2:0]  _EVAL_69,
  input         _EVAL_70,
  input  [1:0]  _EVAL_71,
  output        _EVAL_72,
  output [7:0]  _EVAL_73,
  input  [2:0]  _EVAL_74,
  input         _EVAL_75,
  output [10:0] _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output [2:0]  _EVAL_79,
  output [31:0] _EVAL_80
);
  assign _EVAL_73 = _EVAL_27;
  assign _EVAL_49 = _EVAL_50;
  assign _EVAL = _EVAL_35;
  assign _EVAL_76 = _EVAL_4;
  assign _EVAL_59 = {{1'd0}, _EVAL_23};
  assign _EVAL_26 = _EVAL_37;
  assign _EVAL_57 = _EVAL_46[2:0];
  assign _EVAL_0 = _EVAL_10;
  assign _EVAL_66 = _EVAL_42;
  assign _EVAL_72 = _EVAL_6;
  assign _EVAL_38 = _EVAL_40;
  assign _EVAL_55 = _EVAL_64;
  assign _EVAL_2 = _EVAL_14;
  assign _EVAL_65 = _EVAL_70;
  assign _EVAL_79 = _EVAL_69;
  assign _EVAL_52 = _EVAL_12;
  assign _EVAL_80 = _EVAL_1;
  assign _EVAL_61 = _EVAL_17;
  assign _EVAL_43 = _EVAL_47;
  assign _EVAL_48 = _EVAL_24;
  assign _EVAL_67 = _EVAL_51;
  assign _EVAL_41 = _EVAL_68;
  assign _EVAL_29 = _EVAL_62;
  assign _EVAL_31 = _EVAL_75;
  assign _EVAL_32 = _EVAL_56;
  assign _EVAL_54 = _EVAL_71;
  assign _EVAL_9 = _EVAL_8;
  assign _EVAL_11 = _EVAL_28;
  assign _EVAL_30 = _EVAL_5;
  assign _EVAL_33 = _EVAL_63;
  assign _EVAL_16 = _EVAL_44;
  assign _EVAL_39 = _EVAL_19;
  assign _EVAL_20 = {{1'd0}, _EVAL_74};
  assign _EVAL_7 = _EVAL_36;
  assign _EVAL_3 = _EVAL_21;
  assign _EVAL_13 = _EVAL_60;
  assign _EVAL_78 = _EVAL_25;
  assign _EVAL_45 = _EVAL_15[2:0];
  assign _EVAL_77 = _EVAL_22;
  assign _EVAL_53 = _EVAL_34;
  assign _EVAL_18 = _EVAL_58;
endmodule
