//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_87(
  input         _EVAL,
  input         _EVAL_0,
  input  [63:0] _EVAL_1,
  output        _EVAL_2,
  output [7:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [63:0] _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  output [63:0] _EVAL_15,
  output [2:0]  _EVAL_16,
  output        _EVAL_17,
  input  [2:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  output [2:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input  [7:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  output [2:0]  _EVAL_30,
  output [63:0] _EVAL_31,
  output        _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input  [2:0]  _EVAL_35,
  output [2:0]  _EVAL_36
);
  assign _EVAL_20 = _EVAL_6;
  assign _EVAL_29 = _EVAL_33;
  assign _EVAL_36 = _EVAL_19;
  assign _EVAL_17 = _EVAL;
  assign _EVAL_27 = _EVAL_13;
  assign _EVAL_22 = _EVAL_9;
  assign _EVAL_21 = _EVAL_34;
  assign _EVAL_8 = _EVAL_23;
  assign _EVAL_3 = _EVAL_26;
  assign _EVAL_32 = _EVAL_25;
  assign _EVAL_31 = _EVAL_5;
  assign _EVAL_28 = _EVAL_12;
  assign _EVAL_7 = _EVAL_14;
  assign _EVAL_16 = _EVAL_18;
  assign _EVAL_15 = _EVAL_1;
  assign _EVAL_11 = _EVAL_35;
  assign _EVAL_30 = _EVAL_4;
  assign _EVAL_2 = _EVAL_0;
endmodule
