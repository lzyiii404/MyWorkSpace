//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_169_assert(
  input  [1:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [11:0] _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  input         _EVAL_7,
  input  [11:0] _EVAL_8,
  input  [29:0] _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [3:0]  _EVAL_16
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_19;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_1;
  reg [29:0] _EVAL_50;
  reg [31:0] _RAND_2;
  reg [11:0] _EVAL_59;
  reg [31:0] _RAND_3;
  reg [2335:0] _EVAL_79;
  reg [2335:0] _RAND_4;
  reg  _EVAL_126;
  reg [31:0] _RAND_5;
  reg  _EVAL_135;
  reg [31:0] _RAND_6;
  reg [2:0] _EVAL_160;
  reg [31:0] _RAND_7;
  reg  _EVAL_165;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_175;
  reg [31:0] _RAND_9;
  reg [1:0] _EVAL_194;
  reg [31:0] _RAND_10;
  reg [11:0] _EVAL_204;
  reg [31:0] _RAND_11;
  reg [1:0] _EVAL_231;
  reg [31:0] _RAND_12;
  reg  _EVAL_243;
  reg [31:0] _RAND_13;
  reg [31:0] _EVAL_253;
  reg [31:0] _RAND_14;
  wire [29:0] _EVAL_113;
  wire [30:0] _EVAL_49;
  wire  _EVAL_34;
  wire  _EVAL_222;
  wire  _EVAL_43;
  wire  _EVAL_101;
  wire  _EVAL_91;
  wire  _EVAL_183;
  wire  _EVAL_38;
  wire  _EVAL_221;
  wire  _EVAL_197;
  wire [4095:0] _EVAL_142;
  wire [4095:0] _EVAL_66;
  wire [2335:0] _EVAL_57;
  wire [2335:0] _EVAL_212;
  wire [2335:0] _EVAL_249;
  wire  _EVAL_95;
  wire  _EVAL_90;
  wire  _EVAL_205;
  wire  _EVAL_60;
  wire  _EVAL_230;
  wire  _EVAL_33;
  wire [1:0] _EVAL_24;
  wire [1:0] _EVAL_186;
  wire  _EVAL_224;
  wire  _EVAL_37;
  wire  _EVAL_72;
  wire  _EVAL_55;
  wire  _EVAL_118;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_209;
  wire  _EVAL_139;
  wire  _EVAL_25;
  wire  _EVAL_149;
  wire  _EVAL_77;
  wire  _EVAL_115;
  wire  _EVAL_96;
  wire  _EVAL_56;
  wire  _EVAL_251;
  wire  _EVAL_233;
  wire  _EVAL_89;
  wire  _EVAL_158;
  wire  _EVAL_192;
  wire  _EVAL_114;
  wire  _EVAL_69;
  wire [3:0] _EVAL_23;
  wire  _EVAL_148;
  wire  _EVAL_218;
  wire  _EVAL_80;
  wire  _EVAL_202;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_88;
  wire  _EVAL_107;
  wire  _EVAL_147;
  wire  _EVAL_154;
  wire [4095:0] _EVAL_159;
  wire [4095:0] _EVAL_170;
  wire [2335:0] _EVAL_73;
  wire  _EVAL_220;
  wire  _EVAL_252;
  wire  _EVAL_74;
  wire  _EVAL_157;
  wire  _EVAL_188;
  wire  _EVAL_198;
  wire  _EVAL_61;
  wire  _EVAL_110;
  wire  _EVAL_151;
  wire  _EVAL_123;
  wire  _EVAL_240;
  wire  _EVAL_199;
  wire  _EVAL_239;
  wire  _EVAL_150;
  wire  _EVAL_30;
  wire  _EVAL_168;
  wire  _EVAL_68;
  wire  _EVAL_67;
  wire  _EVAL_161;
  wire  _EVAL_103;
  wire  _EVAL_116;
  wire  _EVAL_195;
  wire  _EVAL_131;
  wire  _EVAL_26;
  wire  _EVAL_119;
  wire [2335:0] _EVAL_121;
  wire  _EVAL_132;
  wire  _EVAL_179;
  wire  _EVAL_18;
  wire  _EVAL_102;
  wire [31:0] _EVAL_85;
  wire [3:0] _EVAL_146;
  wire  _EVAL_20;
  wire  _EVAL_185;
  wire  _EVAL_122;
  wire  _EVAL_181;
  wire  _EVAL_143;
  wire  _EVAL_106;
  wire  _EVAL_117;
  wire  _EVAL_225;
  wire  _EVAL_70;
  wire [4:0] _EVAL_169;
  wire [1:0] _EVAL_93;
  wire [1:0] _EVAL_153;
  wire  _EVAL_206;
  wire  _EVAL_29;
  wire  _EVAL_81;
  wire  _EVAL_200;
  wire  _EVAL_241;
  wire  _EVAL_171;
  wire  _EVAL_104;
  wire  _EVAL_27;
  wire  _EVAL_223;
  wire  _EVAL_144;
  wire  _EVAL_17;
  wire  _EVAL_162;
  wire  _EVAL_207;
  wire  _EVAL_174;
  wire  _EVAL_39;
  wire  _EVAL_219;
  wire  _EVAL_189;
  wire [2335:0] _EVAL_182;
  wire [2335:0] _EVAL_35;
  wire [2335:0] _EVAL_244;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_141;
  wire  _EVAL_105;
  wire  _EVAL_45;
  wire  _EVAL_193;
  wire  _EVAL_138;
  wire  _EVAL_36;
  wire  _EVAL_245;
  wire  _EVAL_42;
  wire  _EVAL_246;
  wire  _EVAL_40;
  wire  _EVAL_125;
  wire  _EVAL_140;
  wire  _EVAL_211;
  wire [29:0] _EVAL_62;
  wire [29:0] _EVAL_226;
  wire  _EVAL_164;
  wire  _EVAL_130;
  wire  _EVAL_127;
  wire  _EVAL_31;
  wire  _EVAL_217;
  wire  _EVAL_247;
  wire  _EVAL_46;
  wire [30:0] _EVAL_203;
  wire [30:0] _EVAL_177;
  wire  _EVAL_134;
  wire  _EVAL_120;
  wire  _EVAL_75;
  wire  _EVAL_109;
  wire  _EVAL_52;
  wire  _EVAL_184;
  wire  _EVAL_98;
  wire  _EVAL_228;
  wire  _EVAL_136;
  wire  _EVAL_133;
  wire  _EVAL_108;
  wire  _EVAL_163;
  wire  _EVAL_99;
  wire  _EVAL_71;
  wire [3:0] _EVAL_44;
  wire [3:0] _EVAL_145;
  wire  _EVAL_236;
  wire  _EVAL_232;
  wire  _EVAL_82;
  wire  _EVAL_227;
  wire  _EVAL_216;
  wire  _EVAL_94;
  wire  _EVAL_210;
  wire  _EVAL_64;
  wire  _EVAL_248;
  wire  _EVAL_180;
  wire  _EVAL_83;
  wire  _EVAL_137;
  wire  _EVAL_214;
  wire  _EVAL_128;
  wire  _EVAL_201;
  wire  _EVAL_87;
  wire  _EVAL_213;
  wire  _EVAL_215;
  wire  _EVAL_63;
  wire  _EVAL_152;
  wire  _EVAL_129;
  wire  _EVAL_41;
  wire  _EVAL_178;
  wire  _EVAL_84;
  wire  _EVAL_176;
  wire  _EVAL_97;
  wire  _EVAL_208;
  wire  _EVAL_54;
  wire  _EVAL_124;
  wire  _EVAL_58;
  wire  _EVAL_112;
  wire  _EVAL_51;
  wire  _EVAL_196;
  wire  _EVAL_78;
  wire  _EVAL_53;
  wire  _EVAL_235;
  wire  _EVAL_173;
  wire  _EVAL_76;
  wire  _EVAL_229;
  wire  _EVAL_86;
  wire  _EVAL_250;
  wire  _EVAL_92;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_113 = _EVAL_9 ^ 30'h20000000;
  assign _EVAL_49 = {1'b0,$signed(_EVAL_113)};
  assign _EVAL_34 = _EVAL_13 & _EVAL_2;
  assign _EVAL_222 = _EVAL_135 == 1'h0;
  assign _EVAL_43 = _EVAL_34 & _EVAL_222;
  assign _EVAL_101 = _EVAL_5 == 1'h0;
  assign _EVAL_91 = _EVAL_101 | _EVAL_10;
  assign _EVAL_183 = _EVAL_91 | _EVAL_3;
  assign _EVAL_38 = _EVAL_183 == 1'h0;
  assign _EVAL_221 = _EVAL_19 == 1'h0;
  assign _EVAL_197 = _EVAL_8 == _EVAL_204;
  assign _EVAL_142 = 4096'h1 << _EVAL_4;
  assign _EVAL_66 = _EVAL_43 ? _EVAL_142 : 4096'h0;
  assign _EVAL_57 = _EVAL_66[2335:0];
  assign _EVAL_212 = _EVAL_57 | _EVAL_79;
  assign _EVAL_249 = _EVAL_212 >> _EVAL_8;
  assign _EVAL_95 = _EVAL_249[0];
  assign _EVAL_90 = _EVAL_15 <= 3'h3;
  assign _EVAL_205 = _EVAL_1 == _EVAL_160;
  assign _EVAL_60 = _EVAL_205 | _EVAL_3;
  assign _EVAL_230 = _EVAL_6 >= 2'h2;
  assign _EVAL_33 = _EVAL_6[0];
  assign _EVAL_24 = 2'h1 << _EVAL_33;
  assign _EVAL_186 = _EVAL_24 | 2'h1;
  assign _EVAL_224 = _EVAL_186[1];
  assign _EVAL_37 = _EVAL_9[1];
  assign _EVAL_72 = _EVAL_224 & _EVAL_37;
  assign _EVAL_55 = _EVAL_230 | _EVAL_72;
  assign _EVAL_118 = _EVAL_186[0];
  assign _EVAL_190 = _EVAL_9[0];
  assign _EVAL_191 = _EVAL_37 & _EVAL_190;
  assign _EVAL_209 = _EVAL_118 & _EVAL_191;
  assign _EVAL_139 = _EVAL_55 | _EVAL_209;
  assign _EVAL_25 = _EVAL_190 == 1'h0;
  assign _EVAL_149 = _EVAL_37 & _EVAL_25;
  assign _EVAL_77 = _EVAL_118 & _EVAL_149;
  assign _EVAL_115 = _EVAL_55 | _EVAL_77;
  assign _EVAL_96 = _EVAL_37 == 1'h0;
  assign _EVAL_56 = _EVAL_224 & _EVAL_96;
  assign _EVAL_251 = _EVAL_230 | _EVAL_56;
  assign _EVAL_233 = _EVAL_96 & _EVAL_190;
  assign _EVAL_89 = _EVAL_118 & _EVAL_233;
  assign _EVAL_158 = _EVAL_251 | _EVAL_89;
  assign _EVAL_192 = _EVAL_96 & _EVAL_25;
  assign _EVAL_114 = _EVAL_118 & _EVAL_192;
  assign _EVAL_69 = _EVAL_251 | _EVAL_114;
  assign _EVAL_23 = {_EVAL_139,_EVAL_115,_EVAL_158,_EVAL_69};
  assign _EVAL_148 = _EVAL_16 == _EVAL_23;
  assign _EVAL_218 = _EVAL_148 | _EVAL_3;
  assign _EVAL_80 = _EVAL_218 == 1'h0;
  assign _EVAL_202 = _EVAL_3 == 1'h0;
  assign _EVAL_237 = _EVAL_7 & _EVAL_11;
  assign _EVAL_238 = _EVAL_165 == 1'h0;
  assign _EVAL_88 = _EVAL_237 & _EVAL_238;
  assign _EVAL_107 = _EVAL_0 == 3'h6;
  assign _EVAL_147 = _EVAL_107 == 1'h0;
  assign _EVAL_154 = _EVAL_88 & _EVAL_147;
  assign _EVAL_159 = 4096'h1 << _EVAL_8;
  assign _EVAL_170 = _EVAL_154 ? _EVAL_159 : 4096'h0;
  assign _EVAL_73 = _EVAL_170[2335:0];
  assign _EVAL_220 = _EVAL_5 == _EVAL_243;
  assign _EVAL_252 = _EVAL_220 | _EVAL_3;
  assign _EVAL_74 = _EVAL_252 == 1'h0;
  assign _EVAL_157 = _EVAL == _EVAL_231;
  assign _EVAL_188 = _EVAL_157 | _EVAL_3;
  assign _EVAL_198 = _EVAL_188 == 1'h0;
  assign _EVAL_61 = _EVAL_57 != 2336'h0;
  assign _EVAL_110 = _EVAL_61 == 1'h0;
  assign _EVAL_151 = _EVAL_165 - 1'h1;
  assign _EVAL_123 = _EVAL_1 == 3'h5;
  assign _EVAL_240 = _EVAL_2 & _EVAL_123;
  assign _EVAL_199 = _EVAL_15 == _EVAL_175;
  assign _EVAL_239 = _EVAL_199 | _EVAL_3;
  assign _EVAL_150 = _EVAL_221 == 1'h0;
  assign _EVAL_30 = _EVAL_2 & _EVAL_150;
  assign _EVAL_168 = _EVAL_0 == 3'h4;
  assign _EVAL_68 = _EVAL_11 & _EVAL_168;
  assign _EVAL_67 = _EVAL_15 <= 3'h4;
  assign _EVAL_161 = _EVAL_67 | _EVAL_3;
  assign _EVAL_103 = _EVAL_161 == 1'h0;
  assign _EVAL_116 = _EVAL_0 == _EVAL_32;
  assign _EVAL_195 = _EVAL_1 == 3'h2;
  assign _EVAL_131 = _EVAL_2 & _EVAL_195;
  assign _EVAL_26 = _EVAL_126 == 1'h0;
  assign _EVAL_119 = _EVAL_126 - 1'h1;
  assign _EVAL_121 = _EVAL_79 >> _EVAL_4;
  assign _EVAL_132 = _EVAL_121[0];
  assign _EVAL_179 = _EVAL_132 == 1'h0;
  assign _EVAL_18 = _EVAL_179 | _EVAL_3;
  assign _EVAL_102 = _EVAL_18 == 1'h0;
  assign _EVAL_85 = _EVAL_253 + 32'h1;
  assign _EVAL_146 = ~ _EVAL_16;
  assign _EVAL_20 = _EVAL_0 == 3'h0;
  assign _EVAL_185 = _EVAL_11 & _EVAL_20;
  assign _EVAL_122 = _EVAL_15 != 3'h0;
  assign _EVAL_181 = _EVAL_122 | _EVAL_3;
  assign _EVAL_143 = _EVAL_181 == 1'h0;
  assign _EVAL_106 = _EVAL_0 <= 3'h6;
  assign _EVAL_117 = _EVAL_15 <= 3'h2;
  assign _EVAL_225 = _EVAL_117 | _EVAL_3;
  assign _EVAL_70 = _EVAL_225 == 1'h0;
  assign _EVAL_169 = 5'h3 << _EVAL_6;
  assign _EVAL_93 = _EVAL_169[1:0];
  assign _EVAL_153 = ~ _EVAL_93;
  assign _EVAL_206 = _EVAL_1 == 3'h7;
  assign _EVAL_29 = _EVAL_2 & _EVAL_206;
  assign _EVAL_81 = _EVAL_79 != 2336'h0;
  assign _EVAL_200 = _EVAL_81 == 1'h0;
  assign _EVAL_241 = plusarg_reader_out == 32'h0;
  assign _EVAL_171 = _EVAL_200 | _EVAL_241;
  assign _EVAL_104 = _EVAL_253 < plusarg_reader_out;
  assign _EVAL_27 = _EVAL_171 | _EVAL_104;
  assign _EVAL_223 = _EVAL_27 | _EVAL_3;
  assign _EVAL_144 = _EVAL_101 | _EVAL_3;
  assign _EVAL_17 = _EVAL_144 == 1'h0;
  assign _EVAL_162 = _EVAL_0 == 3'h5;
  assign _EVAL_207 = _EVAL_4 <= 12'h91f;
  assign _EVAL_174 = _EVAL_26 == 1'h0;
  assign _EVAL_39 = _EVAL_57 != _EVAL_73;
  assign _EVAL_219 = _EVAL_39 | _EVAL_110;
  assign _EVAL_189 = _EVAL_219 | _EVAL_3;
  assign _EVAL_182 = _EVAL_79 | _EVAL_57;
  assign _EVAL_35 = ~ _EVAL_73;
  assign _EVAL_244 = _EVAL_182 & _EVAL_35;
  assign _EVAL_166 = _EVAL_135 - 1'h1;
  assign _EVAL_167 = _EVAL_116 | _EVAL_3;
  assign _EVAL_141 = _EVAL_9 == _EVAL_50;
  assign _EVAL_105 = _EVAL_141 | _EVAL_3;
  assign _EVAL_45 = _EVAL_105 == 1'h0;
  assign _EVAL_193 = _EVAL_6 <= 2'h2;
  assign _EVAL_138 = _EVAL_230 | _EVAL_3;
  assign _EVAL_36 = _EVAL_138 == 1'h0;
  assign _EVAL_245 = _EVAL_1 == 3'h0;
  assign _EVAL_42 = _EVAL_2 & _EVAL_245;
  assign _EVAL_246 = _EVAL_12 == 1'h0;
  assign _EVAL_40 = _EVAL_246 | _EVAL_3;
  assign _EVAL_125 = _EVAL_40 == 1'h0;
  assign _EVAL_140 = _EVAL_6 == _EVAL_194;
  assign _EVAL_211 = _EVAL_140 | _EVAL_3;
  assign _EVAL_62 = {{28'd0}, _EVAL_153};
  assign _EVAL_226 = _EVAL_9 & _EVAL_62;
  assign _EVAL_164 = _EVAL_226 == 30'h0;
  assign _EVAL_130 = _EVAL_164 | _EVAL_3;
  assign _EVAL_127 = _EVAL_130 == 1'h0;
  assign _EVAL_31 = _EVAL_207 | _EVAL_3;
  assign _EVAL_217 = _EVAL_10 == 1'h0;
  assign _EVAL_247 = _EVAL_0 == 3'h1;
  assign _EVAL_46 = _EVAL_11 & _EVAL_247;
  assign _EVAL_203 = $signed(_EVAL_49) & $signed(-31'sh2000);
  assign _EVAL_177 = $signed(_EVAL_203);
  assign _EVAL_134 = $signed(_EVAL_177) == $signed(31'sh0);
  assign _EVAL_120 = _EVAL_193 & _EVAL_134;
  assign _EVAL_75 = _EVAL_120 | _EVAL_3;
  assign _EVAL_109 = _EVAL_75 == 1'h0;
  assign _EVAL_52 = _EVAL_31 == 1'h0;
  assign _EVAL_184 = _EVAL_34 | _EVAL_237;
  assign _EVAL_98 = _EVAL_197 | _EVAL_3;
  assign _EVAL_228 = _EVAL_98 == 1'h0;
  assign _EVAL_136 = _EVAL_60 == 1'h0;
  assign _EVAL_133 = _EVAL >= 2'h2;
  assign _EVAL_108 = _EVAL_133 | _EVAL_3;
  assign _EVAL_163 = _EVAL_108 == 1'h0;
  assign _EVAL_99 = _EVAL_1 == 3'h4;
  assign _EVAL_71 = _EVAL_211 == 1'h0;
  assign _EVAL_44 = ~ _EVAL_23;
  assign _EVAL_145 = _EVAL_16 & _EVAL_44;
  assign _EVAL_236 = _EVAL_223 == 1'h0;
  assign _EVAL_232 = _EVAL_106 | _EVAL_3;
  assign _EVAL_82 = _EVAL_15 == 3'h0;
  assign _EVAL_227 = _EVAL_82 | _EVAL_3;
  assign _EVAL_216 = _EVAL_237 & _EVAL_26;
  assign _EVAL_94 = _EVAL_232 == 1'h0;
  assign _EVAL_210 = _EVAL_2 & _EVAL_99;
  assign _EVAL_64 = _EVAL_217 | _EVAL_3;
  assign _EVAL_248 = _EVAL_64 == 1'h0;
  assign _EVAL_180 = _EVAL_4 == _EVAL_59;
  assign _EVAL_83 = _EVAL_180 | _EVAL_3;
  assign _EVAL_137 = _EVAL_83 == 1'h0;
  assign _EVAL_214 = _EVAL_0 == 3'h2;
  assign _EVAL_128 = _EVAL_11 & _EVAL_214;
  assign _EVAL_201 = _EVAL_145 == 4'h0;
  assign _EVAL_87 = _EVAL_201 | _EVAL_3;
  assign _EVAL_213 = _EVAL_19 - 1'h1;
  assign _EVAL_215 = _EVAL_1 == 3'h1;
  assign _EVAL_63 = _EVAL_239 == 1'h0;
  assign _EVAL_152 = _EVAL_90 | _EVAL_3;
  assign _EVAL_129 = _EVAL_95 | _EVAL_3;
  assign _EVAL_41 = _EVAL_11 & _EVAL_107;
  assign _EVAL_178 = _EVAL_146 == 4'h0;
  assign _EVAL_84 = _EVAL_8 <= 12'h91f;
  assign _EVAL_176 = _EVAL_84 | _EVAL_3;
  assign _EVAL_97 = _EVAL_176 == 1'h0;
  assign _EVAL_208 = _EVAL_1 == 3'h3;
  assign _EVAL_54 = _EVAL_2 & _EVAL_208;
  assign _EVAL_124 = _EVAL_129 == 1'h0;
  assign _EVAL_58 = _EVAL_1 == 3'h6;
  assign _EVAL_112 = _EVAL_2 & _EVAL_58;
  assign _EVAL_51 = _EVAL_87 == 1'h0;
  assign _EVAL_196 = _EVAL_34 & _EVAL_221;
  assign _EVAL_78 = _EVAL_189 == 1'h0;
  assign _EVAL_53 = _EVAL_227 == 1'h0;
  assign _EVAL_235 = _EVAL_2 & _EVAL_215;
  assign _EVAL_173 = _EVAL_167 == 1'h0;
  assign _EVAL_76 = _EVAL_178 | _EVAL_3;
  assign _EVAL_229 = _EVAL_76 == 1'h0;
  assign _EVAL_86 = _EVAL_152 == 1'h0;
  assign _EVAL_250 = _EVAL_11 & _EVAL_162;
  assign _EVAL_92 = _EVAL_11 & _EVAL_174;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_32 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_50 = _RAND_2[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_59 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {73{`RANDOM}};
  _EVAL_79 = _RAND_4[2335:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_126 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_135 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_160 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_165 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_175 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_194 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_204 = _RAND_11[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_231 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_243 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_253 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL_3) begin
      _EVAL_19 <= 1'h0;
    end else begin
      if (_EVAL_34) begin
        if (_EVAL_221) begin
          _EVAL_19 <= 1'h0;
        end else begin
          _EVAL_19 <= _EVAL_213;
        end
      end
    end
    if (_EVAL_216) begin
      _EVAL_32 <= _EVAL_0;
    end
    if (_EVAL_196) begin
      _EVAL_50 <= _EVAL_9;
    end
    if (_EVAL_196) begin
      _EVAL_59 <= _EVAL_4;
    end
    if (_EVAL_3) begin
      _EVAL_79 <= 2336'h0;
    end else begin
      _EVAL_79 <= _EVAL_244;
    end
    if (_EVAL_3) begin
      _EVAL_126 <= 1'h0;
    end else begin
      if (_EVAL_237) begin
        if (_EVAL_26) begin
          _EVAL_126 <= 1'h0;
        end else begin
          _EVAL_126 <= _EVAL_119;
        end
      end
    end
    if (_EVAL_3) begin
      _EVAL_135 <= 1'h0;
    end else begin
      if (_EVAL_34) begin
        if (_EVAL_222) begin
          _EVAL_135 <= 1'h0;
        end else begin
          _EVAL_135 <= _EVAL_166;
        end
      end
    end
    if (_EVAL_196) begin
      _EVAL_160 <= _EVAL_1;
    end
    if (_EVAL_3) begin
      _EVAL_165 <= 1'h0;
    end else begin
      if (_EVAL_237) begin
        if (_EVAL_238) begin
          _EVAL_165 <= 1'h0;
        end else begin
          _EVAL_165 <= _EVAL_151;
        end
      end
    end
    if (_EVAL_196) begin
      _EVAL_175 <= _EVAL_15;
    end
    if (_EVAL_196) begin
      _EVAL_194 <= _EVAL_6;
    end
    if (_EVAL_216) begin
      _EVAL_204 <= _EVAL_8;
    end
    if (_EVAL_216) begin
      _EVAL_231 <= _EVAL;
    end
    if (_EVAL_216) begin
      _EVAL_243 <= _EVAL_5;
    end
    if (_EVAL_3) begin
      _EVAL_253 <= 32'h0;
    end else begin
      if (_EVAL_184) begin
        _EVAL_253 <= 32'h0;
      end else begin
        _EVAL_253 <= _EVAL_85;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f01144e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a1110a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6486ad9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e2338c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab104118)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38e775a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f96225c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b607afc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d9e0d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4abb63a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ada157b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a6d3b0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(305ff33b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80ed0412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f41dbbc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ebd3e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de4efa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6b4229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(712e6f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b62ac05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de0937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec7dc1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e56d81f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16db40b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f8e54cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5973c421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd8beefc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df5ce594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c7cbef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e9bb47c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(852043e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33d13a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c29ce2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75c6894a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79f15155)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(461d4869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28f7b2d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd9f8982)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc6f7efd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b759a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3db41353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(984e3368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928433de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(788dcbf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0f1ad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc9b2a8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a23dce3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f69fe626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6934e7b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(298429ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(764fe0df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c64ea4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4b13773)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7197070)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b619d3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(382bd8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2e71f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a74407f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a9963f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6845e0d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a4f9179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdb425f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f3cccf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cc751f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d66e03f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(319f2bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7cbd3ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c59fc98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3ee7b0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2caa6da2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(128cd404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18aed00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65c12d87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb7bdddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fadacc9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf7b4aea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d2f79c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c52d786)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9401d31d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1df0753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
