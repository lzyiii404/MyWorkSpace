//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_247_assert(
  input  [7:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input  [7:0]  _EVAL_1,
  input  [24:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14
);
  wire [31:0] plusarg_reader_out;
  reg [2:0] _EVAL_16;
  reg [31:0] _RAND_0;
  reg [2:0] _EVAL_36;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_44;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_52;
  reg [31:0] _RAND_3;
  reg [135:0] _EVAL_63;
  reg [159:0] _RAND_4;
  reg [2:0] _EVAL_64;
  reg [31:0] _RAND_5;
  reg [7:0] _EVAL_92;
  reg [31:0] _RAND_6;
  reg [7:0] _EVAL_207;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_239;
  reg [31:0] _RAND_8;
  reg [2:0] _EVAL_242;
  reg [31:0] _RAND_9;
  reg [3:0] _EVAL_250;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_258;
  reg [31:0] _RAND_11;
  reg [3:0] _EVAL_278;
  reg [31:0] _RAND_12;
  reg [24:0] _EVAL_289;
  reg [31:0] _RAND_13;
  wire  _EVAL_147;
  wire  _EVAL_37;
  wire  _EVAL_259;
  wire  _EVAL_165;
  wire  _EVAL_146;
  wire  _EVAL_228;
  wire  _EVAL_287;
  wire [4:0] _EVAL_98;
  wire  _EVAL_96;
  wire [2:0] _EVAL_54;
  wire  _EVAL_80;
  wire  _EVAL_88;
  wire  _EVAL_177;
  wire  _EVAL_298;
  wire  _EVAL_75;
  wire  _EVAL_162;
  wire  _EVAL_172;
  wire  _EVAL_46;
  wire  _EVAL_186;
  wire  _EVAL_45;
  wire  _EVAL_295;
  wire  _EVAL_179;
  wire  _EVAL_142;
  wire  _EVAL_184;
  wire  _EVAL_48;
  wire  _EVAL_27;
  wire  _EVAL_120;
  wire  _EVAL_257;
  wire  _EVAL_280;
  wire  _EVAL_241;
  wire  _EVAL_200;
  wire  _EVAL_91;
  wire  _EVAL_89;
  wire  _EVAL_185;
  wire  _EVAL_18;
  wire  _EVAL_193;
  wire  _EVAL_150;
  wire  _EVAL_132;
  wire [4:0] _EVAL_149;
  wire  _EVAL_153;
  wire [2:0] _EVAL_247;
  wire  _EVAL_222;
  wire  _EVAL_90;
  wire  _EVAL_283;
  wire  _EVAL_156;
  wire  _EVAL_249;
  wire  _EVAL_238;
  wire  _EVAL_190;
  wire  _EVAL_224;
  wire  _EVAL_166;
  wire  _EVAL_231;
  wire  _EVAL_271;
  wire  _EVAL_269;
  wire [12:0] _EVAL_73;
  wire [5:0] _EVAL_17;
  wire [5:0] _EVAL_164;
  wire [135:0] _EVAL_215;
  wire  _EVAL_148;
  wire  _EVAL_124;
  wire  _EVAL_35;
  wire  _EVAL_181;
  wire  _EVAL_266;
  wire [24:0] _EVAL_131;
  wire [25:0] _EVAL_201;
  wire [25:0] _EVAL_274;
  wire [25:0] _EVAL_182;
  wire  _EVAL_110;
  wire  _EVAL_155;
  wire  _EVAL_125;
  wire  _EVAL_67;
  wire  _EVAL_134;
  wire  _EVAL_251;
  wire  _EVAL_236;
  wire [12:0] _EVAL_229;
  wire  _EVAL_101;
  wire  _EVAL_49;
  wire  _EVAL_94;
  wire [3:0] _EVAL_116;
  wire  _EVAL_76;
  wire  _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_296;
  wire  _EVAL_29;
  wire  _EVAL_55;
  wire  _EVAL_303;
  wire  _EVAL_151;
  wire  _EVAL_191;
  wire  _EVAL_135;
  wire  _EVAL_255;
  wire  _EVAL_99;
  wire  _EVAL_38;
  wire [1:0] _EVAL_129;
  wire [1:0] _EVAL_168;
  wire  _EVAL_286;
  wire  _EVAL_87;
  wire  _EVAL_30;
  wire  _EVAL_43;
  wire  _EVAL_62;
  wire  _EVAL_84;
  wire  _EVAL_246;
  wire [5:0] _EVAL_270;
  wire [5:0] _EVAL_93;
  wire  _EVAL_108;
  wire  _EVAL_223;
  wire  _EVAL_139;
  wire  _EVAL_82;
  wire  _EVAL_176;
  wire  _EVAL_42;
  wire  _EVAL_279;
  wire  _EVAL_144;
  wire  _EVAL_103;
  wire  _EVAL_206;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_210;
  wire  _EVAL_192;
  wire  _EVAL_58;
  wire  _EVAL_171;
  wire  _EVAL_232;
  wire  _EVAL_66;
  wire  _EVAL_72;
  wire  _EVAL_77;
  wire  _EVAL_234;
  wire  _EVAL_71;
  wire  _EVAL_272;
  wire  _EVAL_130;
  wire  _EVAL_21;
  wire  _EVAL_152;
  wire  _EVAL_304;
  wire  _EVAL_56;
  wire  _EVAL_197;
  wire  _EVAL_199;
  wire  _EVAL_211;
  wire  _EVAL_187;
  wire  _EVAL_15;
  wire [3:0] _EVAL_145;
  wire [3:0] _EVAL_260;
  wire [3:0] _EVAL_170;
  wire  _EVAL_69;
  wire  _EVAL_34;
  wire  _EVAL_20;
  wire  _EVAL_294;
  wire  _EVAL_198;
  wire [255:0] _EVAL_138;
  wire [255:0] _EVAL_163;
  wire [135:0] _EVAL_154;
  wire [255:0] _EVAL_107;
  wire [255:0] _EVAL_284;
  wire [135:0] _EVAL_212;
  wire  _EVAL_243;
  wire  _EVAL_51;
  wire  _EVAL_180;
  wire  _EVAL_104;
  wire  _EVAL_78;
  wire  _EVAL_262;
  wire  _EVAL_32;
  wire  _EVAL_40;
  wire  _EVAL_106;
  wire  _EVAL_219;
  wire  _EVAL_57;
  wire  _EVAL_221;
  wire [3:0] _EVAL_174;
  wire  _EVAL_118;
  wire  _EVAL_28;
  wire  _EVAL_133;
  wire [135:0] _EVAL_256;
  wire  _EVAL_216;
  wire  _EVAL_204;
  wire  _EVAL_244;
  wire  _EVAL_22;
  wire  _EVAL_175;
  wire  _EVAL_301;
  wire  _EVAL_95;
  wire  _EVAL_275;
  wire  _EVAL_136;
  wire  _EVAL_202;
  wire  _EVAL_209;
  wire  _EVAL_276;
  wire  _EVAL_141;
  wire [135:0] _EVAL_189;
  wire  _EVAL_237;
  wire  _EVAL_268;
  wire [3:0] _EVAL_208;
  wire [24:0] _EVAL_169;
  wire [24:0] _EVAL_288;
  wire  _EVAL_188;
  wire  _EVAL_97;
  wire  _EVAL_79;
  wire  _EVAL_81;
  wire  _EVAL_159;
  wire [3:0] _EVAL_121;
  wire  _EVAL_240;
  wire  _EVAL_161;
  wire  _EVAL_195;
  wire  _EVAL_160;
  wire  _EVAL_158;
  wire  _EVAL_205;
  wire  _EVAL_230;
  wire  _EVAL_263;
  wire  _EVAL_297;
  wire  _EVAL_53;
  wire  _EVAL_194;
  wire  _EVAL_217;
  wire [3:0] _EVAL_50;
  wire [3:0] _EVAL_39;
  wire [135:0] _EVAL_122;
  wire [31:0] _EVAL_83;
  wire [3:0] _EVAL_302;
  wire  _EVAL_167;
  wire  _EVAL_127;
  wire  _EVAL_293;
  wire  _EVAL_261;
  wire  _EVAL_65;
  wire  _EVAL_285;
  wire  _EVAL_85;
  wire [135:0] _EVAL_264;
  wire  _EVAL_299;
  wire  _EVAL_102;
  wire  _EVAL_203;
  wire  _EVAL_47;
  wire  _EVAL_112;
  wire  _EVAL_105;
  wire  _EVAL_128;
  wire  _EVAL_140;
  wire  _EVAL_290;
  wire  _EVAL_277;
  wire  _EVAL_245;
  wire  _EVAL_273;
  wire  _EVAL_74;
  wire [135:0] _EVAL_233;
  wire  _EVAL_143;
  wire  _EVAL_292;
  wire  _EVAL_248;
  wire  _EVAL_213;
  wire  _EVAL_291;
  wire  _EVAL_33;
  wire  _EVAL_126;
  wire  _EVAL_137;
  wire  _EVAL_24;
  wire  _EVAL_226;
  wire  _EVAL_254;
  wire  _EVAL_23;
  wire  _EVAL_114;
  wire  _EVAL_178;
  wire  _EVAL_267;
  wire  _EVAL_265;
  wire  _EVAL_41;
  wire  _EVAL_19;
  wire  _EVAL_252;
  wire  _EVAL_115;
  wire  _EVAL_183;
  wire  _EVAL_86;
  wire  _EVAL_235;
  wire  _EVAL_26;
  wire  _EVAL_282;
  wire  _EVAL_113;
  wire  _EVAL_100;
  wire  _EVAL_119;
  wire  _EVAL_281;
  wire  _EVAL_220;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_147 = _EVAL_10 == _EVAL_64;
  assign _EVAL_37 = _EVAL_147 | _EVAL_3;
  assign _EVAL_259 = _EVAL_12 == 3'h0;
  assign _EVAL_165 = _EVAL_1 == 8'h48;
  assign _EVAL_146 = _EVAL == 8'h48;
  assign _EVAL_228 = _EVAL == 8'h40;
  assign _EVAL_287 = _EVAL_146 | _EVAL_228;
  assign _EVAL_98 = _EVAL[7:3];
  assign _EVAL_96 = _EVAL_98 == 5'h8;
  assign _EVAL_54 = _EVAL[2:0];
  assign _EVAL_80 = 3'h1 <= _EVAL_54;
  assign _EVAL_88 = _EVAL_96 & _EVAL_80;
  assign _EVAL_177 = _EVAL_287 | _EVAL_88;
  assign _EVAL_298 = _EVAL == 8'h20;
  assign _EVAL_75 = _EVAL_177 | _EVAL_298;
  assign _EVAL_162 = _EVAL_98 == 5'h0;
  assign _EVAL_172 = _EVAL_75 | _EVAL_162;
  assign _EVAL_46 = _EVAL_98 == 5'h1;
  assign _EVAL_186 = _EVAL_172 | _EVAL_46;
  assign _EVAL_45 = _EVAL_98 == 5'h2;
  assign _EVAL_295 = _EVAL_186 | _EVAL_45;
  assign _EVAL_179 = _EVAL_98 == 5'h3;
  assign _EVAL_142 = _EVAL_295 | _EVAL_179;
  assign _EVAL_184 = _EVAL == 8'h80;
  assign _EVAL_48 = _EVAL_142 | _EVAL_184;
  assign _EVAL_27 = _EVAL_98 == 5'h10;
  assign _EVAL_120 = _EVAL_27 & _EVAL_80;
  assign _EVAL_257 = _EVAL_48 | _EVAL_120;
  assign _EVAL_280 = _EVAL_257 | _EVAL_3;
  assign _EVAL_241 = _EVAL_280 == 1'h0;
  assign _EVAL_200 = _EVAL_4 & _EVAL_11;
  assign _EVAL_91 = _EVAL_250 == 4'h0;
  assign _EVAL_89 = _EVAL_200 & _EVAL_91;
  assign _EVAL_185 = _EVAL_12 == 3'h6;
  assign _EVAL_18 = _EVAL_185 == 1'h0;
  assign _EVAL_193 = _EVAL_89 & _EVAL_18;
  assign _EVAL_150 = _EVAL_1 == 8'h40;
  assign _EVAL_132 = _EVAL_165 | _EVAL_150;
  assign _EVAL_149 = _EVAL_1[7:3];
  assign _EVAL_153 = _EVAL_149 == 5'h8;
  assign _EVAL_247 = _EVAL_1[2:0];
  assign _EVAL_222 = 3'h1 <= _EVAL_247;
  assign _EVAL_90 = _EVAL_153 & _EVAL_222;
  assign _EVAL_283 = _EVAL_132 | _EVAL_90;
  assign _EVAL_156 = _EVAL_1 == 8'h20;
  assign _EVAL_249 = _EVAL_283 | _EVAL_156;
  assign _EVAL_238 = _EVAL_149 == 5'h0;
  assign _EVAL_190 = _EVAL_249 | _EVAL_238;
  assign _EVAL_224 = _EVAL_149 == 5'h1;
  assign _EVAL_166 = _EVAL_190 | _EVAL_224;
  assign _EVAL_231 = _EVAL_278 == 4'h0;
  assign _EVAL_271 = _EVAL_231 == 1'h0;
  assign _EVAL_269 = _EVAL_9 & _EVAL_271;
  assign _EVAL_73 = 13'h3f << _EVAL_5;
  assign _EVAL_17 = _EVAL_73[5:0];
  assign _EVAL_164 = ~ _EVAL_17;
  assign _EVAL_215 = _EVAL_63 >> _EVAL;
  assign _EVAL_148 = _EVAL_215[0];
  assign _EVAL_124 = _EVAL_10 != 3'h0;
  assign _EVAL_35 = _EVAL_124 | _EVAL_3;
  assign _EVAL_181 = _EVAL_35 == 1'h0;
  assign _EVAL_266 = _EVAL_11 & _EVAL_185;
  assign _EVAL_131 = _EVAL_2 ^ 25'h1900000;
  assign _EVAL_201 = {1'b0,$signed(_EVAL_131)};
  assign _EVAL_274 = $signed(_EVAL_201) & $signed(-26'sh2000);
  assign _EVAL_182 = $signed(_EVAL_274);
  assign _EVAL_110 = _EVAL_63 != 136'h0;
  assign _EVAL_155 = _EVAL_110 == 1'h0;
  assign _EVAL_125 = plusarg_reader_out == 32'h0;
  assign _EVAL_67 = _EVAL_155 | _EVAL_125;
  assign _EVAL_134 = _EVAL_52 < plusarg_reader_out;
  assign _EVAL_251 = _EVAL_67 | _EVAL_134;
  assign _EVAL_236 = _EVAL_251 | _EVAL_3;
  assign _EVAL_229 = 13'h3f << _EVAL_0;
  assign _EVAL_101 = _EVAL_10 <= 3'h2;
  assign _EVAL_49 = _EVAL_101 | _EVAL_3;
  assign _EVAL_94 = _EVAL_49 == 1'h0;
  assign _EVAL_116 = ~ _EVAL_13;
  assign _EVAL_76 = _EVAL_116 == 4'h0;
  assign _EVAL_68 = _EVAL_76 | _EVAL_3;
  assign _EVAL_70 = _EVAL_68 == 1'h0;
  assign _EVAL_296 = _EVAL_6 == 3'h4;
  assign _EVAL_29 = _EVAL_9 & _EVAL_296;
  assign _EVAL_55 = _EVAL_8 & _EVAL_9;
  assign _EVAL_303 = _EVAL_55 | _EVAL_200;
  assign _EVAL_151 = _EVAL_2[1];
  assign _EVAL_191 = _EVAL_151 == 1'h0;
  assign _EVAL_135 = _EVAL_2[0];
  assign _EVAL_255 = _EVAL_135 == 1'h0;
  assign _EVAL_99 = _EVAL_191 & _EVAL_255;
  assign _EVAL_38 = _EVAL_5[0];
  assign _EVAL_129 = 2'h1 << _EVAL_38;
  assign _EVAL_168 = _EVAL_129 | 2'h1;
  assign _EVAL_286 = _EVAL_168[1];
  assign _EVAL_87 = _EVAL_5 >= 3'h2;
  assign _EVAL_30 = _EVAL_0 == _EVAL_258;
  assign _EVAL_43 = _EVAL_149 == 5'h2;
  assign _EVAL_62 = _EVAL_166 | _EVAL_43;
  assign _EVAL_84 = _EVAL_149 == 5'h3;
  assign _EVAL_246 = _EVAL_62 | _EVAL_84;
  assign _EVAL_270 = _EVAL_229[5:0];
  assign _EVAL_93 = ~ _EVAL_270;
  assign _EVAL_108 = _EVAL_12 == 3'h1;
  assign _EVAL_223 = _EVAL_11 & _EVAL_108;
  assign _EVAL_139 = 3'h6 == _EVAL_5;
  assign _EVAL_82 = _EVAL_228 ? _EVAL_139 : 1'h0;
  assign _EVAL_176 = _EVAL_184 ? _EVAL_139 : 1'h0;
  assign _EVAL_42 = _EVAL_82 | _EVAL_176;
  assign _EVAL_279 = _EVAL_168[0];
  assign _EVAL_144 = _EVAL_151 & _EVAL_135;
  assign _EVAL_103 = _EVAL_279 & _EVAL_144;
  assign _EVAL_206 = _EVAL_5 == _EVAL_16;
  assign _EVAL_60 = _EVAL_206 | _EVAL_3;
  assign _EVAL_61 = _EVAL_60 == 1'h0;
  assign _EVAL_210 = _EVAL_3 == 1'h0;
  assign _EVAL_192 = _EVAL_286 & _EVAL_191;
  assign _EVAL_58 = _EVAL_87 | _EVAL_192;
  assign _EVAL_171 = _EVAL_279 & _EVAL_99;
  assign _EVAL_232 = _EVAL_58 | _EVAL_171;
  assign _EVAL_66 = _EVAL_11 & _EVAL_259;
  assign _EVAL_72 = _EVAL_12 == 3'h5;
  assign _EVAL_77 = _EVAL_6 == 3'h7;
  assign _EVAL_234 = _EVAL_9 & _EVAL_77;
  assign _EVAL_71 = _EVAL_6 == 3'h2;
  assign _EVAL_272 = _EVAL_9 & _EVAL_71;
  assign _EVAL_130 = _EVAL_10 == 3'h0;
  assign _EVAL_21 = _EVAL_286 & _EVAL_151;
  assign _EVAL_152 = _EVAL_87 | _EVAL_21;
  assign _EVAL_304 = _EVAL_152 | _EVAL_103;
  assign _EVAL_56 = _EVAL_151 & _EVAL_255;
  assign _EVAL_197 = _EVAL_279 & _EVAL_56;
  assign _EVAL_199 = _EVAL_152 | _EVAL_197;
  assign _EVAL_211 = _EVAL_191 & _EVAL_135;
  assign _EVAL_187 = _EVAL_279 & _EVAL_211;
  assign _EVAL_15 = _EVAL_58 | _EVAL_187;
  assign _EVAL_145 = {_EVAL_304,_EVAL_199,_EVAL_15,_EVAL_232};
  assign _EVAL_260 = ~ _EVAL_145;
  assign _EVAL_170 = _EVAL_13 & _EVAL_260;
  assign _EVAL_69 = _EVAL_170 == 4'h0;
  assign _EVAL_34 = _EVAL_69 | _EVAL_3;
  assign _EVAL_20 = _EVAL_34 == 1'h0;
  assign _EVAL_294 = _EVAL_239 == 4'h0;
  assign _EVAL_198 = _EVAL_55 & _EVAL_294;
  assign _EVAL_138 = 256'h1 << _EVAL;
  assign _EVAL_163 = _EVAL_198 ? _EVAL_138 : 256'h0;
  assign _EVAL_154 = _EVAL_163[135:0];
  assign _EVAL_107 = 256'h1 << _EVAL_1;
  assign _EVAL_284 = _EVAL_193 ? _EVAL_107 : 256'h0;
  assign _EVAL_212 = _EVAL_284[135:0];
  assign _EVAL_243 = _EVAL_154 != _EVAL_212;
  assign _EVAL_51 = _EVAL_154 != 136'h0;
  assign _EVAL_180 = _EVAL_51 == 1'h0;
  assign _EVAL_104 = _EVAL_243 | _EVAL_180;
  assign _EVAL_78 = _EVAL_104 | _EVAL_3;
  assign _EVAL_262 = _EVAL_12 == 3'h2;
  assign _EVAL_32 = _EVAL_1 == 8'h80;
  assign _EVAL_40 = _EVAL_246 | _EVAL_32;
  assign _EVAL_106 = _EVAL_149 == 5'h10;
  assign _EVAL_219 = _EVAL_106 & _EVAL_222;
  assign _EVAL_57 = _EVAL_40 | _EVAL_219;
  assign _EVAL_221 = _EVAL_6[2];
  assign _EVAL_174 = _EVAL_44 - 4'h1;
  assign _EVAL_118 = _EVAL_7 == 1'h0;
  assign _EVAL_28 = _EVAL_118 | _EVAL_3;
  assign _EVAL_133 = _EVAL_28 == 1'h0;
  assign _EVAL_256 = ~ _EVAL_212;
  assign _EVAL_216 = _EVAL_13 == _EVAL_145;
  assign _EVAL_204 = _EVAL_216 | _EVAL_3;
  assign _EVAL_244 = _EVAL_204 == 1'h0;
  assign _EVAL_22 = _EVAL_0 >= 3'h2;
  assign _EVAL_175 = _EVAL_5 <= 3'h2;
  assign _EVAL_301 = $signed(_EVAL_182) == $signed(26'sh0);
  assign _EVAL_95 = _EVAL_175 & _EVAL_301;
  assign _EVAL_275 = _EVAL_95 | _EVAL_3;
  assign _EVAL_136 = _EVAL_30 | _EVAL_3;
  assign _EVAL_202 = _EVAL_136 == 1'h0;
  assign _EVAL_209 = _EVAL_148 == 1'h0;
  assign _EVAL_276 = _EVAL_209 | _EVAL_3;
  assign _EVAL_141 = _EVAL_276 == 1'h0;
  assign _EVAL_189 = _EVAL_154 | _EVAL_63;
  assign _EVAL_237 = _EVAL_44 == 4'h0;
  assign _EVAL_268 = _EVAL_12[0];
  assign _EVAL_208 = _EVAL_93[5:2];
  assign _EVAL_169 = {{19'd0}, _EVAL_164};
  assign _EVAL_288 = _EVAL_2 & _EVAL_169;
  assign _EVAL_188 = _EVAL_288 == 25'h0;
  assign _EVAL_97 = _EVAL_275 == 1'h0;
  assign _EVAL_79 = _EVAL_10 <= 3'h3;
  assign _EVAL_81 = _EVAL_79 | _EVAL_3;
  assign _EVAL_159 = _EVAL_81 == 1'h0;
  assign _EVAL_121 = _EVAL_250 - 4'h1;
  assign _EVAL_240 = _EVAL_2 == _EVAL_289;
  assign _EVAL_161 = _EVAL_240 | _EVAL_3;
  assign _EVAL_195 = _EVAL_12 <= 3'h6;
  assign _EVAL_160 = _EVAL_195 | _EVAL_3;
  assign _EVAL_158 = _EVAL_6 == 3'h0;
  assign _EVAL_205 = _EVAL_9 & _EVAL_158;
  assign _EVAL_230 = _EVAL_6 == 3'h3;
  assign _EVAL_263 = _EVAL_57 | _EVAL_3;
  assign _EVAL_297 = _EVAL_263 == 1'h0;
  assign _EVAL_53 = _EVAL_12 == 3'h4;
  assign _EVAL_194 = _EVAL_11 & _EVAL_53;
  assign _EVAL_217 = _EVAL_221 == 1'h0;
  assign _EVAL_50 = _EVAL_164[5:2];
  assign _EVAL_39 = _EVAL_239 - 4'h1;
  assign _EVAL_122 = _EVAL_63 | _EVAL_154;
  assign _EVAL_83 = _EVAL_52 + 32'h1;
  assign _EVAL_302 = _EVAL_278 - 4'h1;
  assign _EVAL_167 = _EVAL_10 <= 3'h4;
  assign _EVAL_127 = _EVAL_167 | _EVAL_3;
  assign _EVAL_293 = _EVAL_9 & _EVAL_230;
  assign _EVAL_261 = _EVAL_161 == 1'h0;
  assign _EVAL_65 = _EVAL_1 == _EVAL_207;
  assign _EVAL_285 = _EVAL_65 | _EVAL_3;
  assign _EVAL_85 = _EVAL == _EVAL_92;
  assign _EVAL_264 = _EVAL_189 >> _EVAL_1;
  assign _EVAL_299 = _EVAL_264[0];
  assign _EVAL_102 = _EVAL_285 == 1'h0;
  assign _EVAL_203 = _EVAL_6 == 3'h6;
  assign _EVAL_47 = _EVAL_78 == 1'h0;
  assign _EVAL_112 = _EVAL_42 | _EVAL_3;
  assign _EVAL_105 = _EVAL_12 == _EVAL_36;
  assign _EVAL_128 = _EVAL_105 | _EVAL_3;
  assign _EVAL_140 = _EVAL_128 == 1'h0;
  assign _EVAL_290 = _EVAL_5 <= 3'h6;
  assign _EVAL_277 = _EVAL_112 == 1'h0;
  assign _EVAL_245 = _EVAL_87 | _EVAL_3;
  assign _EVAL_273 = _EVAL_245 == 1'h0;
  assign _EVAL_74 = _EVAL_200 & _EVAL_237;
  assign _EVAL_233 = _EVAL_122 & _EVAL_256;
  assign _EVAL_143 = _EVAL_237 == 1'h0;
  assign _EVAL_292 = _EVAL_11 & _EVAL_143;
  assign _EVAL_248 = _EVAL_11 & _EVAL_72;
  assign _EVAL_213 = _EVAL_6 == 3'h5;
  assign _EVAL_291 = _EVAL_9 & _EVAL_213;
  assign _EVAL_33 = _EVAL_85 | _EVAL_3;
  assign _EVAL_126 = _EVAL_33 == 1'h0;
  assign _EVAL_137 = _EVAL_22 | _EVAL_3;
  assign _EVAL_24 = _EVAL_6 == 3'h1;
  assign _EVAL_226 = _EVAL_9 & _EVAL_24;
  assign _EVAL_254 = _EVAL_137 == 1'h0;
  assign _EVAL_23 = _EVAL_6 == _EVAL_242;
  assign _EVAL_114 = _EVAL_23 | _EVAL_3;
  assign _EVAL_178 = _EVAL_114 == 1'h0;
  assign _EVAL_267 = _EVAL_299 | _EVAL_3;
  assign _EVAL_265 = _EVAL_267 == 1'h0;
  assign _EVAL_41 = _EVAL_37 == 1'h0;
  assign _EVAL_19 = _EVAL_55 & _EVAL_231;
  assign _EVAL_252 = _EVAL_188 | _EVAL_3;
  assign _EVAL_115 = _EVAL_130 | _EVAL_3;
  assign _EVAL_183 = _EVAL_115 == 1'h0;
  assign _EVAL_86 = _EVAL_290 & _EVAL_301;
  assign _EVAL_235 = _EVAL_127 == 1'h0;
  assign _EVAL_26 = _EVAL_252 == 1'h0;
  assign _EVAL_282 = _EVAL_86 | _EVAL_3;
  assign _EVAL_113 = _EVAL_236 == 1'h0;
  assign _EVAL_100 = _EVAL_9 & _EVAL_203;
  assign _EVAL_119 = _EVAL_160 == 1'h0;
  assign _EVAL_281 = _EVAL_282 == 1'h0;
  assign _EVAL_220 = _EVAL_11 & _EVAL_262;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_16 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_36 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_44 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_52 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {5{`RANDOM}};
  _EVAL_63 = _RAND_4[135:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_64 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_92 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_207 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_239 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_242 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_250 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_258 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_278 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_289 = _RAND_13[24:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_14) begin
    if (_EVAL_19) begin
      _EVAL_16 <= _EVAL_5;
    end
    if (_EVAL_74) begin
      _EVAL_36 <= _EVAL_12;
    end
    if (_EVAL_3) begin
      _EVAL_44 <= 4'h0;
    end else begin
      if (_EVAL_200) begin
        if (_EVAL_237) begin
          if (_EVAL_268) begin
            _EVAL_44 <= _EVAL_208;
          end else begin
            _EVAL_44 <= 4'h0;
          end
        end else begin
          _EVAL_44 <= _EVAL_174;
        end
      end
    end
    if (_EVAL_3) begin
      _EVAL_52 <= 32'h0;
    end else begin
      if (_EVAL_303) begin
        _EVAL_52 <= 32'h0;
      end else begin
        _EVAL_52 <= _EVAL_83;
      end
    end
    if (_EVAL_3) begin
      _EVAL_63 <= 136'h0;
    end else begin
      _EVAL_63 <= _EVAL_233;
    end
    if (_EVAL_19) begin
      _EVAL_64 <= _EVAL_10;
    end
    if (_EVAL_19) begin
      _EVAL_92 <= _EVAL;
    end
    if (_EVAL_74) begin
      _EVAL_207 <= _EVAL_1;
    end
    if (_EVAL_3) begin
      _EVAL_239 <= 4'h0;
    end else begin
      if (_EVAL_55) begin
        if (_EVAL_294) begin
          if (_EVAL_217) begin
            _EVAL_239 <= _EVAL_50;
          end else begin
            _EVAL_239 <= 4'h0;
          end
        end else begin
          _EVAL_239 <= _EVAL_39;
        end
      end
    end
    if (_EVAL_19) begin
      _EVAL_242 <= _EVAL_6;
    end
    if (_EVAL_3) begin
      _EVAL_250 <= 4'h0;
    end else begin
      if (_EVAL_200) begin
        if (_EVAL_91) begin
          if (_EVAL_268) begin
            _EVAL_250 <= _EVAL_208;
          end else begin
            _EVAL_250 <= 4'h0;
          end
        end else begin
          _EVAL_250 <= _EVAL_121;
        end
      end
    end
    if (_EVAL_74) begin
      _EVAL_258 <= _EVAL_0;
    end
    if (_EVAL_3) begin
      _EVAL_278 <= 4'h0;
    end else begin
      if (_EVAL_55) begin
        if (_EVAL_231) begin
          if (_EVAL_217) begin
            _EVAL_278 <= _EVAL_50;
          end else begin
            _EVAL_278 <= 4'h0;
          end
        end else begin
          _EVAL_278 <= _EVAL_302;
        end
      end
    end
    if (_EVAL_19) begin
      _EVAL_289 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d73dc71b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8359307f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d064cb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb466fd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afd2c886)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd56365)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31549671)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9709458)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d500830)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58f6b63d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f4b273e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90e74cf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7711bde8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca35c8df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0acd675)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee2e798c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2444e67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c21e302)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aafb825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96f22b7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8569c97b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20cb536f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(806c47a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e84580ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33a04dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e44834e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60035d5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da80cc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4459a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fa546d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4ffabb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63140195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8062f310)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6073644b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14c307ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3918b28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b53ce7bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfdc534d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6e395b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4557d22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc8ddaeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60312637)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39927b0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38775631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(723b7e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bca910f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b24c00d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3850cfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(785716ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e54727a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a35074d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2fd5be9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac11c63e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78fddb5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6772f24f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(667e5af0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16efb9fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(458d2fec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2120db8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92118c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6c8b41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c981a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6f05cc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94c3eac8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1614927c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5191b543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(309e6c64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c11e3844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7830b8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55514007)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eebf182c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(968b4802)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
