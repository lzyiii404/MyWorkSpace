//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive__EVAL_191_assert(
  input        _EVAL,
  input        _EVAL_0,
  input  [2:0] _EVAL_1,
  input  [2:0] _EVAL_2,
  input        _EVAL_3,
  input  [3:0] _EVAL_4,
  input  [6:0] _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8
);
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_12;
  reg [31:0] _RAND_0;
  reg [6:0] _EVAL_30;
  reg [31:0] _RAND_1;
  reg  _EVAL_43;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_48;
  reg [31:0] _RAND_3;
  reg  _EVAL_61;
  reg [31:0] _RAND_4;
  reg [2:0] _EVAL_95;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_103;
  reg [31:0] _RAND_6;
  reg  _EVAL_105;
  reg [31:0] _RAND_7;
  reg  _EVAL_107;
  reg [31:0] _RAND_8;
  wire  _EVAL_104;
  wire  _EVAL_37;
  wire  _EVAL_108;
  wire  _EVAL_15;
  wire [6:0] _EVAL_79;
  wire  _EVAL_72;
  wire  _EVAL_120;
  wire  _EVAL_77;
  wire  _EVAL_55;
  wire  _EVAL_32;
  wire  _EVAL_25;
  wire  _EVAL_27;
  wire [1:0] _EVAL_57;
  wire  _EVAL_111;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_49;
  wire  _EVAL_16;
  wire  _EVAL_75;
  wire  _EVAL_65;
  wire  _EVAL_82;
  wire [1:0] _EVAL_31;
  wire  _EVAL_51;
  wire  _EVAL_46;
  wire  _EVAL_129;
  wire  _EVAL_22;
  wire  _EVAL_66;
  wire  _EVAL_87;
  wire  _EVAL_53;
  wire [6:0] _EVAL_24;
  wire [7:0] _EVAL_117;
  wire [7:0] _EVAL_115;
  wire [7:0] _EVAL_18;
  wire  _EVAL_78;
  wire [6:0] _EVAL_67;
  wire [7:0] _EVAL_76;
  wire [7:0] _EVAL_36;
  wire [7:0] _EVAL_29;
  wire  _EVAL_123;
  wire  _EVAL_63;
  wire  _EVAL_39;
  wire  _EVAL_21;
  wire  _EVAL_42;
  wire  _EVAL_74;
  wire  _EVAL_35;
  wire  _EVAL_17;
  wire  _EVAL_90;
  wire  _EVAL_89;
  wire  _EVAL_38;
  wire [31:0] _EVAL_126;
  wire  _EVAL_93;
  wire  _EVAL_52;
  wire  _EVAL_62;
  wire  _EVAL_50;
  wire  _EVAL_97;
  wire  _EVAL_125;
  wire  _EVAL_19;
  wire  _EVAL_60;
  wire [3:0] _EVAL_81;
  wire  _EVAL_73;
  wire  _EVAL_99;
  wire  _EVAL_128;
  wire  _EVAL_98;
  wire  _EVAL_118;
  wire  _EVAL_59;
  wire  _EVAL_121;
  wire  _EVAL_80;
  wire  _EVAL_127;
  wire  _EVAL_102;
  wire  _EVAL_45;
  wire  _EVAL_56;
  wire  _EVAL_116;
  wire  _EVAL_122;
  wire  _EVAL_34;
  wire  _EVAL_40;
  wire  _EVAL_14;
  wire  _EVAL_114;
  wire  _EVAL_47;
  wire  _EVAL_100;
  wire  _EVAL_96;
  wire  _EVAL_64;
  wire  _EVAL_130;
  wire  _EVAL_44;
  wire  _EVAL_83;
  wire  _EVAL_23;
  wire  _EVAL_119;
  wire  _EVAL_91;
  wire  _EVAL_94;
  wire  _EVAL_71;
  wire  _EVAL_54;
  wire  _EVAL_26;
  wire  _EVAL_70;
  wire  _EVAL_11;
  wire  _EVAL_33;
  wire  _EVAL_69;
  wire  _EVAL_84;
  wire  _EVAL_10;
  wire  _EVAL_112;
  wire  _EVAL_101;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_104 = _EVAL_1 == _EVAL_95;
  assign _EVAL_37 = _EVAL_104 | _EVAL;
  assign _EVAL_108 = _EVAL_1 == 3'h2;
  assign _EVAL_15 = _EVAL_1 == 3'h4;
  assign _EVAL_79 = _EVAL_5 & 7'h3;
  assign _EVAL_72 = _EVAL_79 == 7'h0;
  assign _EVAL_120 = _EVAL_72 | _EVAL;
  assign _EVAL_77 = _EVAL_5 == _EVAL_30;
  assign _EVAL_55 = _EVAL_77 | _EVAL;
  assign _EVAL_32 = _EVAL_3 & _EVAL_8;
  assign _EVAL_25 = _EVAL_12 == 1'h0;
  assign _EVAL_27 = _EVAL_32 & _EVAL_25;
  assign _EVAL_57 = _EVAL_27 ? 2'h1 : 2'h0;
  assign _EVAL_111 = _EVAL_57[0];
  assign _EVAL_85 = _EVAL_61 | _EVAL_111;
  assign _EVAL_86 = _EVAL_7 & _EVAL_6;
  assign _EVAL_49 = _EVAL_43 == 1'h0;
  assign _EVAL_16 = _EVAL_86 & _EVAL_49;
  assign _EVAL_75 = _EVAL_2 == 3'h6;
  assign _EVAL_65 = _EVAL_75 == 1'h0;
  assign _EVAL_82 = _EVAL_16 & _EVAL_65;
  assign _EVAL_31 = _EVAL_82 ? 2'h1 : 2'h0;
  assign _EVAL_51 = _EVAL_31[0];
  assign _EVAL_46 = ~ _EVAL_51;
  assign _EVAL_129 = _EVAL_85 & _EVAL_46;
  assign _EVAL_22 = _EVAL_105 == 1'h0;
  assign _EVAL_66 = _EVAL_105 - 1'h1;
  assign _EVAL_87 = _EVAL_107 == 1'h0;
  assign _EVAL_53 = _EVAL_107 - 1'h1;
  assign _EVAL_24 = _EVAL_5 ^ 7'h40;
  assign _EVAL_117 = {1'b0,$signed(_EVAL_24)};
  assign _EVAL_115 = $signed(_EVAL_117) & $signed(-8'sh14);
  assign _EVAL_18 = $signed(_EVAL_115);
  assign _EVAL_78 = $signed(_EVAL_18) == $signed(8'sh0);
  assign _EVAL_67 = _EVAL_5 ^ 7'h54;
  assign _EVAL_76 = {1'b0,$signed(_EVAL_67)};
  assign _EVAL_36 = $signed(_EVAL_76) & $signed(-8'sh4);
  assign _EVAL_29 = $signed(_EVAL_36);
  assign _EVAL_123 = $signed(_EVAL_29) == $signed(8'sh0);
  assign _EVAL_63 = _EVAL_78 | _EVAL_123;
  assign _EVAL_39 = _EVAL_63 | _EVAL;
  assign _EVAL_21 = _EVAL_12 - 1'h1;
  assign _EVAL_42 = _EVAL_8 & _EVAL_108;
  assign _EVAL_74 = _EVAL_1 == 3'h0;
  assign _EVAL_35 = _EVAL_1 == 3'h7;
  assign _EVAL_17 = _EVAL_111 | _EVAL_61;
  assign _EVAL_90 = _EVAL_17 | _EVAL;
  assign _EVAL_89 = _EVAL_90 == 1'h0;
  assign _EVAL_38 = _EVAL_87 == 1'h0;
  assign _EVAL_126 = _EVAL_48 + 32'h1;
  assign _EVAL_93 = _EVAL_32 | _EVAL_86;
  assign _EVAL_52 = _EVAL_2 == _EVAL_103;
  assign _EVAL_62 = _EVAL_1 == 3'h3;
  assign _EVAL_50 = _EVAL_8 & _EVAL_62;
  assign _EVAL_97 = _EVAL_8 & _EVAL_15;
  assign _EVAL_125 = _EVAL_1 == 3'h5;
  assign _EVAL_19 = _EVAL_8 & _EVAL_125;
  assign _EVAL_60 = _EVAL_86 & _EVAL_87;
  assign _EVAL_81 = ~ _EVAL_4;
  assign _EVAL_73 = _EVAL_81 == 4'h0;
  assign _EVAL_99 = _EVAL_48 < plusarg_reader_out;
  assign _EVAL_128 = _EVAL_52 | _EVAL;
  assign _EVAL_98 = _EVAL_128 == 1'h0;
  assign _EVAL_118 = _EVAL_61 == 1'h0;
  assign _EVAL_59 = _EVAL_118 | _EVAL;
  assign _EVAL_121 = _EVAL_2 == 3'h5;
  assign _EVAL_80 = _EVAL_43 - 1'h1;
  assign _EVAL_127 = _EVAL_55 == 1'h0;
  assign _EVAL_102 = _EVAL_2 <= 3'h6;
  assign _EVAL_45 = _EVAL_102 | _EVAL;
  assign _EVAL_56 = _EVAL_2 == 3'h4;
  assign _EVAL_116 = _EVAL_73 | _EVAL;
  assign _EVAL_122 = _EVAL_116 == 1'h0;
  assign _EVAL_34 = _EVAL_1 == 3'h1;
  assign _EVAL_40 = _EVAL_8 & _EVAL_74;
  assign _EVAL_14 = _EVAL_22 == 1'h0;
  assign _EVAL_114 = _EVAL_6 & _EVAL_121;
  assign _EVAL_47 = plusarg_reader_out == 32'h0;
  assign _EVAL_100 = _EVAL_118 | _EVAL_47;
  assign _EVAL_96 = _EVAL_4 == 4'hf;
  assign _EVAL_64 = _EVAL_96 | _EVAL;
  assign _EVAL_130 = _EVAL_64 == 1'h0;
  assign _EVAL_44 = _EVAL == 1'h0;
  assign _EVAL_83 = _EVAL_39 == 1'h0;
  assign _EVAL_23 = _EVAL_100 | _EVAL_99;
  assign _EVAL_119 = _EVAL_23 | _EVAL;
  assign _EVAL_91 = _EVAL_119 == 1'h0;
  assign _EVAL_94 = _EVAL_6 & _EVAL_38;
  assign _EVAL_71 = _EVAL_8 & _EVAL_34;
  assign _EVAL_54 = _EVAL_8 & _EVAL_35;
  assign _EVAL_26 = _EVAL_37 == 1'h0;
  assign _EVAL_70 = _EVAL_8 & _EVAL_14;
  assign _EVAL_11 = _EVAL_120 == 1'h0;
  assign _EVAL_33 = _EVAL_1 == 3'h6;
  assign _EVAL_69 = _EVAL_45 == 1'h0;
  assign _EVAL_84 = _EVAL_59 == 1'h0;
  assign _EVAL_10 = _EVAL_6 & _EVAL_56;
  assign _EVAL_112 = _EVAL_32 & _EVAL_22;
  assign _EVAL_101 = _EVAL_8 & _EVAL_33;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_12 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_30 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_43 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_48 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_61 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_95 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_103 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_105 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_107 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_0) begin
    if (_EVAL) begin
      _EVAL_12 <= 1'h0;
    end else begin
      if (_EVAL_32) begin
        if (_EVAL_25) begin
          _EVAL_12 <= 1'h0;
        end else begin
          _EVAL_12 <= _EVAL_21;
        end
      end
    end
    if (_EVAL_112) begin
      _EVAL_30 <= _EVAL_5;
    end
    if (_EVAL) begin
      _EVAL_43 <= 1'h0;
    end else begin
      if (_EVAL_86) begin
        if (_EVAL_49) begin
          _EVAL_43 <= 1'h0;
        end else begin
          _EVAL_43 <= _EVAL_80;
        end
      end
    end
    if (_EVAL) begin
      _EVAL_48 <= 32'h0;
    end else begin
      if (_EVAL_93) begin
        _EVAL_48 <= 32'h0;
      end else begin
        _EVAL_48 <= _EVAL_126;
      end
    end
    if (_EVAL) begin
      _EVAL_61 <= 1'h0;
    end else begin
      _EVAL_61 <= _EVAL_129;
    end
    if (_EVAL_112) begin
      _EVAL_95 <= _EVAL_1;
    end
    if (_EVAL_60) begin
      _EVAL_103 <= _EVAL_2;
    end
    if (_EVAL) begin
      _EVAL_105 <= 1'h0;
    end else begin
      if (_EVAL_32) begin
        if (_EVAL_22) begin
          _EVAL_105 <= 1'h0;
        end else begin
          _EVAL_105 <= _EVAL_66;
        end
      end
    end
    if (_EVAL) begin
      _EVAL_107 <= 1'h0;
    end else begin
      if (_EVAL_86) begin
        if (_EVAL_87) begin
          _EVAL_107 <= 1'h0;
        end else begin
          _EVAL_107 <= _EVAL_53;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0cc5de9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1ed45e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92a1dfd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ce8495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fed8fc1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc37a65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41840a24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e0f3518)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe3ebfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd8ac41a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fac240fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46f47d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6960c2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0df3b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4e62568)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb0ee0c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e10630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b545ca7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62580a4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6023828f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aeb0489)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b55b74d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(137ea209)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d74a700d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_11) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50233e29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b4be3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e94a3e0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d41f7dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed466af0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d00bbce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab6ae77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24475c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b95e39d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74fdaa07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_11) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfc2d21c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
