//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_33(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  output        _EVAL_1,
  output        _EVAL_2,
  output [7:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  output [1:0]  _EVAL_5,
  output [3:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  output [6:0]  _EVAL_12,
  input         _EVAL_13,
  output [2:0]  _EVAL_14,
  input         _EVAL_15,
  input  [1:0]  _EVAL_16,
  output [3:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  output [3:0]  _EVAL_20,
  output [30:0] _EVAL_21,
  input  [10:0] _EVAL_22,
  input  [2:0]  _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  output [31:0] _EVAL_26,
  input         _EVAL_27,
  output        _EVAL_28,
  output [10:0] _EVAL_29,
  output [7:0]  _EVAL_30,
  output        _EVAL_31,
  input  [31:0] _EVAL_32,
  output [2:0]  _EVAL_33,
  input         _EVAL_34,
  output [31:0] _EVAL_35,
  output [2:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  input  [31:0] _EVAL_38,
  input  [2:0]  _EVAL_39,
  output        _EVAL_40,
  input  [6:0]  _EVAL_41,
  output [3:0]  _EVAL_42,
  input  [30:0] _EVAL_43,
  output [3:0]  _EVAL_44,
  output [2:0]  _EVAL_45,
  output [2:0]  _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49,
  output        _EVAL_50,
  input  [10:0] _EVAL_51,
  output [1:0]  _EVAL_52,
  output        _EVAL_53,
  input         _EVAL_54,
  output [30:0] _EVAL_55,
  output [10:0] _EVAL_56,
  output [2:0]  _EVAL_57,
  input  [2:0]  _EVAL_58,
  input         _EVAL_59
);
  wire  Queue__EVAL;
  wire  Queue__EVAL_0;
  wire [3:0] Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire [31:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire [3:0] Queue__EVAL_8;
  wire  Queue__EVAL_9;
  wire [31:0] Queue__EVAL_10;
  wire [10:0] Queue_1__EVAL;
  wire [30:0] Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire [7:0] Queue_1__EVAL_2;
  wire [3:0] Queue_1__EVAL_3;
  wire [1:0] Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire [7:0] Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire [2:0] Queue_1__EVAL_8;
  wire  Queue_1__EVAL_9;
  wire  Queue_1__EVAL_10;
  wire [10:0] Queue_1__EVAL_11;
  wire [30:0] Queue_1__EVAL_12;
  wire  Queue_1__EVAL_13;
  wire [3:0] Queue_1__EVAL_14;
  wire [2:0] Queue_1__EVAL_15;
  wire [2:0] Queue_1__EVAL_16;
  wire [2:0] Queue_1__EVAL_17;
  wire  Queue_1__EVAL_18;
  wire  Queue_1__EVAL_19;
  wire  Queue_1__EVAL_20;
  wire [2:0] Queue_1__EVAL_21;
  reg  _EVAL_89;
  reg [31:0] _RAND_0;
  reg  _EVAL_103;
  reg [31:0] _RAND_1;
  reg [3:0] _EVAL_128;
  reg [31:0] _RAND_2;
  reg  _EVAL_148;
  reg [31:0] _RAND_3;
  reg [3:0] _EVAL_158;
  reg [31:0] _RAND_4;
  reg  _EVAL_196;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_209;
  reg [31:0] _RAND_6;
  reg  _EVAL_212;
  reg [31:0] _RAND_7;
  reg [3:0] _EVAL_252;
  reg [31:0] _RAND_8;
  reg [3:0] _EVAL_286;
  reg [31:0] _RAND_9;
  reg  _EVAL_299;
  reg [31:0] _RAND_10;
  reg  _EVAL_309;
  reg [31:0] _RAND_11;
  reg  _EVAL_314;
  reg [31:0] _RAND_12;
  reg  _EVAL_364;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_377;
  reg [31:0] _RAND_14;
  reg  _EVAL_398;
  reg [31:0] _RAND_15;
  reg  _EVAL_426;
  reg [31:0] _RAND_16;
  reg  _EVAL_430;
  reg [31:0] _RAND_17;
  wire [2:0] _EVAL_166;
  wire [2:0] _EVAL_387;
  wire [2:0] _EVAL_120;
  wire [2:0] _EVAL_350;
  wire [2:0] _EVAL_292;
  wire [2:0] _EVAL_324;
  wire [2:0] _EVAL_359;
  wire [2:0] _EVAL_332;
  wire [2:0] _EVAL_144;
  wire [2:0] _EVAL_64;
  wire [2:0] _EVAL_229;
  wire [2:0] _EVAL_274;
  wire [2:0] _EVAL_291;
  wire [2:0] _EVAL_72;
  wire [2:0] _EVAL_225;
  wire [2:0] _EVAL_242;
  wire [2:0] _EVAL_270;
  wire [2:0] _EVAL_105;
  wire [2:0] _EVAL_337;
  wire [2:0] _EVAL_298;
  wire [2:0] _EVAL_305;
  wire [2:0] _EVAL_78;
  wire [2:0] _EVAL_457;
  wire [2:0] _EVAL_161;
  wire [2:0] _EVAL_369;
  wire [2:0] _EVAL_190;
  wire [2:0] _EVAL_131;
  wire [2:0] _EVAL_422;
  wire [2:0] _EVAL_340;
  wire [2:0] _EVAL_373;
  wire [2:0] _EVAL_94;
  wire [2:0] _EVAL_109;
  wire [2:0] _EVAL_261;
  wire [2:0] _EVAL_421;
  wire [2:0] _EVAL_119;
  wire [2:0] _EVAL_378;
  wire [2:0] _EVAL_362;
  wire [2:0] _EVAL_317;
  wire [2:0] _EVAL_338;
  wire [2:0] _EVAL_189;
  wire [2:0] _EVAL_222;
  wire [2:0] _EVAL_435;
  wire [2:0] _EVAL_344;
  wire [2:0] _EVAL_135;
  wire [2:0] _EVAL_321;
  wire [2:0] _EVAL_442;
  wire [2:0] _EVAL_101;
  wire [2:0] _EVAL_117;
  wire [2:0] _EVAL_112;
  wire [2:0] _EVAL_182;
  wire [2:0] _EVAL_355;
  wire [2:0] _EVAL_175;
  wire [2:0] _EVAL_126;
  wire [2:0] _EVAL_178;
  wire [2:0] _EVAL_456;
  wire [2:0] _EVAL_414;
  wire [2:0] _EVAL_187;
  wire [2:0] _EVAL_444;
  wire [2:0] _EVAL_454;
  wire [2:0] _EVAL_310;
  wire [2:0] _EVAL_287;
  wire [2:0] _EVAL_440;
  wire [2:0] _EVAL_450;
  wire [2:0] _EVAL_184;
  wire [2:0] _EVAL_163;
  wire [7:0] _EVAL_386;
  wire  _EVAL_165;
  wire  _EVAL_403;
  wire  _EVAL_91;
  wire  _EVAL_434;
  wire  _EVAL_315;
  wire  _EVAL_330;
  wire  _EVAL_74;
  wire  _EVAL_308;
  wire  _EVAL_419;
  wire  _EVAL_259;
  wire  _EVAL_154;
  wire  _EVAL_143;
  wire  _EVAL_99;
  wire  _EVAL_409;
  wire  _EVAL_418;
  wire  _EVAL_234;
  wire  _EVAL_250;
  wire  _EVAL_118;
  wire  _EVAL_138;
  wire  _EVAL_416;
  wire  _EVAL_71;
  wire  _EVAL_459;
  wire  _EVAL_179;
  wire  _EVAL_341;
  wire  _EVAL_200;
  wire  _EVAL_280;
  wire  _EVAL_316;
  wire  _EVAL_216;
  wire  _EVAL_235;
  wire  _EVAL_402;
  wire  _EVAL_162;
  wire  _EVAL_153;
  wire  _EVAL_97;
  wire  _EVAL_90;
  wire  _EVAL_169;
  wire  _EVAL_295;
  wire  _EVAL_345;
  wire  _EVAL_436;
  wire  _EVAL_288;
  wire  _EVAL_284;
  wire  _EVAL_157;
  wire  _EVAL_215;
  wire  _EVAL_346;
  wire  _EVAL_336;
  wire  _EVAL_268;
  wire  _EVAL_428;
  wire  _EVAL_382;
  wire  _EVAL_342;
  wire  _EVAL_273;
  wire  _EVAL_420;
  wire  _EVAL_335;
  wire  _EVAL_413;
  wire  _EVAL_352;
  wire  _EVAL_172;
  wire  _EVAL_145;
  wire  _EVAL_220;
  wire  _EVAL_380;
  wire  _EVAL_365;
  wire  _EVAL_255;
  wire  _EVAL_66;
  wire  _EVAL_396;
  wire  _EVAL_63;
  wire  _EVAL_183;
  wire  _EVAL_401;
  wire  _EVAL_443;
  wire  _EVAL_370;
  wire  _EVAL_137;
  wire  _EVAL_264;
  wire  _EVAL_406;
  wire  _EVAL_399;
  wire  _EVAL_244;
  wire  _EVAL_113;
  wire  _EVAL_339;
  wire  _EVAL_69;
  wire  _EVAL_168;
  wire  _EVAL_301;
  wire  _EVAL_447;
  wire  _EVAL_239;
  wire  _EVAL_397;
  wire  _EVAL_203;
  wire  _EVAL_371;
  wire  _EVAL_170;
  wire  _EVAL_210;
  wire  _EVAL_290;
  wire  _EVAL_391;
  wire  _EVAL_226;
  wire  _EVAL_445;
  wire  _EVAL_320;
  wire  _EVAL_151;
  wire  _EVAL_281;
  wire  _EVAL_93;
  wire  _EVAL_171;
  wire  _EVAL_124;
  wire  _EVAL_441;
  wire  _EVAL_347;
  wire  _EVAL_116;
  wire  _EVAL_379;
  wire  _EVAL_205;
  wire  _EVAL_433;
  wire  _EVAL_331;
  wire  _EVAL_155;
  wire  _EVAL_267;
  wire  _EVAL_141;
  wire  _EVAL_455;
  wire  _EVAL_279;
  wire  _EVAL_211;
  wire  _EVAL_123;
  wire  _EVAL_446;
  wire  _EVAL_73;
  wire  _EVAL_388;
  wire  _EVAL_177;
  wire  _EVAL_333;
  wire [2:0] _EVAL_328;
  wire [7:0] _EVAL_204;
  wire  _EVAL_82;
  wire  _EVAL_395;
  wire  _EVAL_424;
  wire  _EVAL_307;
  wire  _EVAL_240;
  wire  _EVAL_429;
  wire  _EVAL_410;
  wire  _EVAL_87;
  wire [3:0] _EVAL_302;
  wire  _EVAL_353;
  wire  _EVAL_110;
  wire  _EVAL_329;
  wire  _EVAL_129;
  wire  _EVAL_88;
  wire  _EVAL_408;
  wire  _EVAL_81;
  wire  _EVAL_458;
  wire  _EVAL_253;
  wire [3:0] _EVAL_357;
  wire  _EVAL_390;
  wire  _EVAL_243;
  wire  _EVAL_407;
  wire  _EVAL_415;
  wire  _EVAL_108;
  wire  _EVAL_263;
  wire  _EVAL_293;
  wire [12:0] _EVAL_366;
  wire  _EVAL_283;
  wire  _EVAL_360;
  wire  _EVAL_160;
  wire  _EVAL_294;
  wire  _EVAL_139;
  wire  _EVAL_351;
  wire  _EVAL_191;
  wire  _EVAL_439;
  wire [9:0] _EVAL_275;
  wire  _EVAL_111;
  wire  _EVAL_152;
  wire [3:0] _EVAL_133;
  wire  _EVAL_206;
  wire [5:0] _EVAL_254;
  wire [5:0] _EVAL_393;
  wire [3:0] _EVAL_62;
  wire [3:0] _EVAL_76;
  wire  _EVAL_136;
  wire  _EVAL_146;
  wire  _EVAL_251;
  wire  _EVAL_334;
  wire  _EVAL_181;
  wire  _EVAL_227;
  wire [6:0] _EVAL_277;
  wire [3:0] _EVAL_276;
  wire [3:0] _EVAL_303;
  wire  _EVAL_202;
  wire  _EVAL_134;
  wire  _EVAL_77;
  wire  _EVAL_392;
  wire  _EVAL_278;
  wire [3:0] _EVAL_199;
  wire  _EVAL_385;
  wire  _EVAL_449;
  wire  _EVAL_404;
  wire  _EVAL_349;
  wire  _EVAL_289;
  wire [3:0] _EVAL_313;
  wire [3:0] _EVAL_356;
  wire [3:0] _EVAL_384;
  wire  _EVAL_300;
  wire  _EVAL_322;
  wire [3:0] _EVAL_311;
  wire [3:0] _EVAL_296;
  wire [16:0] _EVAL_121;
  wire [9:0] _EVAL_282;
  wire [9:0] _EVAL_83;
  wire [9:0] _EVAL_223;
  wire [9:0] _EVAL_100;
  wire  _EVAL_241;
  wire  _EVAL_400;
  wire [3:0] _EVAL_180;
  wire [3:0] _EVAL_427;
  wire [3:0] _EVAL_236;
  wire [2:0] _EVAL_95;
  wire [2:0] _EVAL_431;
  wire [2:0] _EVAL_394;
  wire [2:0] _EVAL_232;
  wire  _EVAL_70;
  wire  _EVAL_192;
  wire  _EVAL_247;
  wire  _EVAL_327;
  wire  _EVAL_319;
  wire [2:0] _EVAL_208;
  wire  _EVAL_147;
  wire [3:0] _EVAL_92;
  wire  _EVAL_285;
  wire [6:0] _EVAL_389;
  wire  _EVAL_306;
  wire  _EVAL_423;
  wire [3:0] _EVAL_85;
  wire [2:0] _EVAL_79;
  wire  _EVAL_194;
  wire  _EVAL_185;
  wire  _EVAL_86;
  wire [3:0] _EVAL_201;
  wire  _EVAL_448;
  SiFive__EVAL_31 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10)
  );
  SiFive__EVAL_32 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14),
    ._EVAL_15(Queue_1__EVAL_15),
    ._EVAL_16(Queue_1__EVAL_16),
    ._EVAL_17(Queue_1__EVAL_17),
    ._EVAL_18(Queue_1__EVAL_18),
    ._EVAL_19(Queue_1__EVAL_19),
    ._EVAL_20(Queue_1__EVAL_20),
    ._EVAL_21(Queue_1__EVAL_21)
  );
  assign _EVAL_166 = 7'h8 == _EVAL_41 ? 3'h4 : 3'h3;
  assign _EVAL_387 = 7'h9 == _EVAL_41 ? 3'h4 : _EVAL_166;
  assign _EVAL_120 = 7'ha == _EVAL_41 ? 3'h4 : _EVAL_387;
  assign _EVAL_350 = 7'hb == _EVAL_41 ? 3'h4 : _EVAL_120;
  assign _EVAL_292 = 7'hc == _EVAL_41 ? 3'h4 : _EVAL_350;
  assign _EVAL_324 = 7'hd == _EVAL_41 ? 3'h4 : _EVAL_292;
  assign _EVAL_359 = 7'he == _EVAL_41 ? 3'h4 : _EVAL_324;
  assign _EVAL_332 = 7'hf == _EVAL_41 ? 3'h4 : _EVAL_359;
  assign _EVAL_144 = 7'h10 == _EVAL_41 ? 3'h5 : _EVAL_332;
  assign _EVAL_64 = 7'h11 == _EVAL_41 ? 3'h5 : _EVAL_144;
  assign _EVAL_229 = 7'h12 == _EVAL_41 ? 3'h5 : _EVAL_64;
  assign _EVAL_274 = 7'h13 == _EVAL_41 ? 3'h5 : _EVAL_229;
  assign _EVAL_291 = 7'h14 == _EVAL_41 ? 3'h5 : _EVAL_274;
  assign _EVAL_72 = 7'h15 == _EVAL_41 ? 3'h5 : _EVAL_291;
  assign _EVAL_225 = 7'h16 == _EVAL_41 ? 3'h5 : _EVAL_72;
  assign _EVAL_242 = 7'h17 == _EVAL_41 ? 3'h5 : _EVAL_225;
  assign _EVAL_270 = 7'h18 == _EVAL_41 ? 3'h6 : _EVAL_242;
  assign _EVAL_105 = 7'h19 == _EVAL_41 ? 3'h6 : _EVAL_270;
  assign _EVAL_337 = 7'h1a == _EVAL_41 ? 3'h6 : _EVAL_105;
  assign _EVAL_298 = 7'h1b == _EVAL_41 ? 3'h6 : _EVAL_337;
  assign _EVAL_305 = 7'h1c == _EVAL_41 ? 3'h6 : _EVAL_298;
  assign _EVAL_78 = 7'h1d == _EVAL_41 ? 3'h6 : _EVAL_305;
  assign _EVAL_457 = 7'h1e == _EVAL_41 ? 3'h6 : _EVAL_78;
  assign _EVAL_161 = 7'h1f == _EVAL_41 ? 3'h6 : _EVAL_457;
  assign _EVAL_369 = 7'h20 == _EVAL_41 ? 3'h1 : _EVAL_161;
  assign _EVAL_190 = 7'h21 == _EVAL_41 ? 3'h0 : _EVAL_369;
  assign _EVAL_131 = 7'h22 == _EVAL_41 ? 3'h0 : _EVAL_190;
  assign _EVAL_422 = 7'h23 == _EVAL_41 ? 3'h0 : _EVAL_131;
  assign _EVAL_340 = 7'h24 == _EVAL_41 ? 3'h0 : _EVAL_422;
  assign _EVAL_373 = 7'h25 == _EVAL_41 ? 3'h0 : _EVAL_340;
  assign _EVAL_94 = 7'h26 == _EVAL_41 ? 3'h0 : _EVAL_373;
  assign _EVAL_109 = 7'h27 == _EVAL_41 ? 3'h0 : _EVAL_94;
  assign _EVAL_261 = 7'h28 == _EVAL_41 ? 3'h0 : _EVAL_109;
  assign _EVAL_421 = 7'h29 == _EVAL_41 ? 3'h0 : _EVAL_261;
  assign _EVAL_119 = 7'h2a == _EVAL_41 ? 3'h0 : _EVAL_421;
  assign _EVAL_378 = 7'h2b == _EVAL_41 ? 3'h0 : _EVAL_119;
  assign _EVAL_362 = 7'h2c == _EVAL_41 ? 3'h0 : _EVAL_378;
  assign _EVAL_317 = 7'h2d == _EVAL_41 ? 3'h0 : _EVAL_362;
  assign _EVAL_338 = 7'h2e == _EVAL_41 ? 3'h0 : _EVAL_317;
  assign _EVAL_189 = 7'h2f == _EVAL_41 ? 3'h0 : _EVAL_338;
  assign _EVAL_222 = 7'h30 == _EVAL_41 ? 3'h0 : _EVAL_189;
  assign _EVAL_435 = 7'h31 == _EVAL_41 ? 3'h0 : _EVAL_222;
  assign _EVAL_344 = 7'h32 == _EVAL_41 ? 3'h0 : _EVAL_435;
  assign _EVAL_135 = 7'h33 == _EVAL_41 ? 3'h0 : _EVAL_344;
  assign _EVAL_321 = 7'h34 == _EVAL_41 ? 3'h0 : _EVAL_135;
  assign _EVAL_442 = 7'h35 == _EVAL_41 ? 3'h0 : _EVAL_321;
  assign _EVAL_101 = 7'h36 == _EVAL_41 ? 3'h0 : _EVAL_442;
  assign _EVAL_117 = 7'h37 == _EVAL_41 ? 3'h0 : _EVAL_101;
  assign _EVAL_112 = 7'h38 == _EVAL_41 ? 3'h0 : _EVAL_117;
  assign _EVAL_182 = 7'h39 == _EVAL_41 ? 3'h0 : _EVAL_112;
  assign _EVAL_355 = 7'h3a == _EVAL_41 ? 3'h0 : _EVAL_182;
  assign _EVAL_175 = 7'h3b == _EVAL_41 ? 3'h0 : _EVAL_355;
  assign _EVAL_126 = 7'h3c == _EVAL_41 ? 3'h0 : _EVAL_175;
  assign _EVAL_178 = 7'h3d == _EVAL_41 ? 3'h0 : _EVAL_126;
  assign _EVAL_456 = 7'h3e == _EVAL_41 ? 3'h0 : _EVAL_178;
  assign _EVAL_414 = 7'h3f == _EVAL_41 ? 3'h0 : _EVAL_456;
  assign _EVAL_187 = 7'h40 == _EVAL_41 ? 3'h7 : _EVAL_414;
  assign _EVAL_444 = 7'h41 == _EVAL_41 ? 3'h2 : _EVAL_187;
  assign _EVAL_454 = 7'h42 == _EVAL_41 ? 3'h2 : _EVAL_444;
  assign _EVAL_310 = 7'h43 == _EVAL_41 ? 3'h2 : _EVAL_454;
  assign _EVAL_287 = 7'h44 == _EVAL_41 ? 3'h2 : _EVAL_310;
  assign _EVAL_440 = 7'h45 == _EVAL_41 ? 3'h2 : _EVAL_287;
  assign _EVAL_450 = 7'h46 == _EVAL_41 ? 3'h2 : _EVAL_440;
  assign _EVAL_184 = 7'h47 == _EVAL_41 ? 3'h2 : _EVAL_450;
  assign _EVAL_163 = 7'h48 == _EVAL_41 ? 3'h0 : _EVAL_184;
  assign _EVAL_386 = 8'h1 << _EVAL_163;
  assign _EVAL_165 = _EVAL_386[0];
  assign _EVAL_403 = _EVAL_377 == 4'h0;
  assign _EVAL_91 = _EVAL_403 == 1'h0;
  assign _EVAL_434 = _EVAL_39[2];
  assign _EVAL_315 = _EVAL_434 == 1'h0;
  assign _EVAL_330 = _EVAL_398 != _EVAL_315;
  assign _EVAL_74 = _EVAL_91 & _EVAL_330;
  assign _EVAL_308 = _EVAL_377 == 4'h8;
  assign _EVAL_419 = _EVAL_74 | _EVAL_308;
  assign _EVAL_259 = _EVAL_252 == 4'h0;
  assign _EVAL_154 = _EVAL_259 == 1'h0;
  assign _EVAL_143 = _EVAL_148 != _EVAL_315;
  assign _EVAL_99 = _EVAL_154 & _EVAL_143;
  assign _EVAL_409 = _EVAL_252 == 4'h8;
  assign _EVAL_418 = _EVAL_99 | _EVAL_409;
  assign _EVAL_234 = _EVAL_158 == 4'h0;
  assign _EVAL_250 = _EVAL_234 == 1'h0;
  assign _EVAL_118 = _EVAL_196 != _EVAL_315;
  assign _EVAL_138 = _EVAL_250 & _EVAL_118;
  assign _EVAL_416 = _EVAL_158 == 4'h8;
  assign _EVAL_71 = _EVAL_138 | _EVAL_416;
  assign _EVAL_459 = _EVAL_128 == 4'h0;
  assign _EVAL_179 = _EVAL_459 == 1'h0;
  assign _EVAL_341 = _EVAL_430 != _EVAL_315;
  assign _EVAL_200 = _EVAL_179 & _EVAL_341;
  assign _EVAL_280 = _EVAL_128 == 4'h8;
  assign _EVAL_316 = _EVAL_200 | _EVAL_280;
  assign _EVAL_216 = 7'h8 == _EVAL_41 ? _EVAL_71 : _EVAL_316;
  assign _EVAL_235 = 7'h9 == _EVAL_41 ? _EVAL_71 : _EVAL_216;
  assign _EVAL_402 = 7'ha == _EVAL_41 ? _EVAL_71 : _EVAL_235;
  assign _EVAL_162 = 7'hb == _EVAL_41 ? _EVAL_71 : _EVAL_402;
  assign _EVAL_153 = 7'hc == _EVAL_41 ? _EVAL_71 : _EVAL_162;
  assign _EVAL_97 = 7'hd == _EVAL_41 ? _EVAL_71 : _EVAL_153;
  assign _EVAL_90 = 7'he == _EVAL_41 ? _EVAL_71 : _EVAL_97;
  assign _EVAL_169 = 7'hf == _EVAL_41 ? _EVAL_71 : _EVAL_90;
  assign _EVAL_295 = 7'h10 == _EVAL_41 ? _EVAL_418 : _EVAL_169;
  assign _EVAL_345 = 7'h11 == _EVAL_41 ? _EVAL_418 : _EVAL_295;
  assign _EVAL_436 = 7'h12 == _EVAL_41 ? _EVAL_418 : _EVAL_345;
  assign _EVAL_288 = 7'h13 == _EVAL_41 ? _EVAL_418 : _EVAL_436;
  assign _EVAL_284 = 7'h14 == _EVAL_41 ? _EVAL_418 : _EVAL_288;
  assign _EVAL_157 = 7'h15 == _EVAL_41 ? _EVAL_418 : _EVAL_284;
  assign _EVAL_215 = 7'h16 == _EVAL_41 ? _EVAL_418 : _EVAL_157;
  assign _EVAL_346 = 7'h17 == _EVAL_41 ? _EVAL_418 : _EVAL_215;
  assign _EVAL_336 = 7'h18 == _EVAL_41 ? _EVAL_419 : _EVAL_346;
  assign _EVAL_268 = 7'h19 == _EVAL_41 ? _EVAL_419 : _EVAL_336;
  assign _EVAL_428 = 7'h1a == _EVAL_41 ? _EVAL_419 : _EVAL_268;
  assign _EVAL_382 = 7'h1b == _EVAL_41 ? _EVAL_419 : _EVAL_428;
  assign _EVAL_342 = 7'h1c == _EVAL_41 ? _EVAL_419 : _EVAL_382;
  assign _EVAL_273 = 7'h1d == _EVAL_41 ? _EVAL_419 : _EVAL_342;
  assign _EVAL_420 = 7'h1e == _EVAL_41 ? _EVAL_419 : _EVAL_273;
  assign _EVAL_335 = 7'h1f == _EVAL_41 ? _EVAL_419 : _EVAL_420;
  assign _EVAL_413 = 7'h20 == _EVAL_41 ? _EVAL_299 : _EVAL_335;
  assign _EVAL_352 = 7'h21 == _EVAL_41 ? 1'h0 : _EVAL_413;
  assign _EVAL_172 = 7'h22 == _EVAL_41 ? 1'h0 : _EVAL_352;
  assign _EVAL_145 = _EVAL_386[6];
  assign _EVAL_220 = Queue_1__EVAL_1;
  assign _EVAL_380 = _EVAL_209 == 3'h0;
  assign _EVAL_365 = _EVAL_380 == 1'h0;
  assign _EVAL_255 = _EVAL_89 != _EVAL_315;
  assign _EVAL_66 = _EVAL_365 & _EVAL_255;
  assign _EVAL_396 = _EVAL_209 == 3'h7;
  assign _EVAL_63 = _EVAL_66 | _EVAL_396;
  assign _EVAL_183 = 7'h23 == _EVAL_41 ? 1'h0 : _EVAL_172;
  assign _EVAL_401 = 7'h24 == _EVAL_41 ? 1'h0 : _EVAL_183;
  assign _EVAL_443 = 7'h25 == _EVAL_41 ? 1'h0 : _EVAL_401;
  assign _EVAL_370 = 7'h26 == _EVAL_41 ? 1'h0 : _EVAL_443;
  assign _EVAL_137 = 7'h27 == _EVAL_41 ? 1'h0 : _EVAL_370;
  assign _EVAL_264 = 7'h28 == _EVAL_41 ? 1'h0 : _EVAL_137;
  assign _EVAL_406 = 7'h29 == _EVAL_41 ? 1'h0 : _EVAL_264;
  assign _EVAL_399 = 7'h2a == _EVAL_41 ? 1'h0 : _EVAL_406;
  assign _EVAL_244 = 7'h2b == _EVAL_41 ? 1'h0 : _EVAL_399;
  assign _EVAL_113 = 7'h2c == _EVAL_41 ? 1'h0 : _EVAL_244;
  assign _EVAL_339 = 7'h2d == _EVAL_41 ? 1'h0 : _EVAL_113;
  assign _EVAL_69 = 7'h2e == _EVAL_41 ? 1'h0 : _EVAL_339;
  assign _EVAL_168 = 7'h2f == _EVAL_41 ? 1'h0 : _EVAL_69;
  assign _EVAL_301 = 7'h30 == _EVAL_41 ? 1'h0 : _EVAL_168;
  assign _EVAL_447 = 7'h31 == _EVAL_41 ? 1'h0 : _EVAL_301;
  assign _EVAL_239 = 7'h32 == _EVAL_41 ? 1'h0 : _EVAL_447;
  assign _EVAL_397 = 7'h33 == _EVAL_41 ? 1'h0 : _EVAL_239;
  assign _EVAL_203 = 7'h34 == _EVAL_41 ? 1'h0 : _EVAL_397;
  assign _EVAL_371 = 7'h35 == _EVAL_41 ? 1'h0 : _EVAL_203;
  assign _EVAL_170 = 7'h36 == _EVAL_41 ? 1'h0 : _EVAL_371;
  assign _EVAL_210 = 7'h37 == _EVAL_41 ? 1'h0 : _EVAL_170;
  assign _EVAL_290 = 7'h38 == _EVAL_41 ? 1'h0 : _EVAL_210;
  assign _EVAL_391 = 7'h39 == _EVAL_41 ? 1'h0 : _EVAL_290;
  assign _EVAL_226 = 7'h3a == _EVAL_41 ? 1'h0 : _EVAL_391;
  assign _EVAL_445 = 7'h3b == _EVAL_41 ? 1'h0 : _EVAL_226;
  assign _EVAL_320 = 7'h3c == _EVAL_41 ? 1'h0 : _EVAL_445;
  assign _EVAL_151 = 7'h3d == _EVAL_41 ? 1'h0 : _EVAL_320;
  assign _EVAL_281 = 7'h3e == _EVAL_41 ? 1'h0 : _EVAL_151;
  assign _EVAL_93 = 7'h3f == _EVAL_41 ? 1'h0 : _EVAL_281;
  assign _EVAL_171 = 7'h40 == _EVAL_41 ? _EVAL_103 : _EVAL_93;
  assign _EVAL_124 = 7'h41 == _EVAL_41 ? _EVAL_63 : _EVAL_171;
  assign _EVAL_441 = 7'h42 == _EVAL_41 ? _EVAL_63 : _EVAL_124;
  assign _EVAL_347 = 7'h43 == _EVAL_41 ? _EVAL_63 : _EVAL_441;
  assign _EVAL_116 = 7'h44 == _EVAL_41 ? _EVAL_63 : _EVAL_347;
  assign _EVAL_379 = 7'h45 == _EVAL_41 ? _EVAL_63 : _EVAL_116;
  assign _EVAL_205 = 7'h46 == _EVAL_41 ? _EVAL_63 : _EVAL_379;
  assign _EVAL_433 = 7'h47 == _EVAL_41 ? _EVAL_63 : _EVAL_205;
  assign _EVAL_331 = 7'h48 == _EVAL_41 ? _EVAL_212 : _EVAL_433;
  assign _EVAL_155 = _EVAL_286 == 4'h0;
  assign _EVAL_267 = _EVAL_331 & _EVAL_155;
  assign _EVAL_141 = _EVAL_267 == 1'h0;
  assign _EVAL_455 = _EVAL_141 & _EVAL_34;
  assign _EVAL_279 = _EVAL_364 == 1'h0;
  assign _EVAL_211 = Queue__EVAL_6;
  assign _EVAL_123 = _EVAL_279 & _EVAL_211;
  assign _EVAL_446 = _EVAL_315 ? _EVAL_123 : 1'h1;
  assign _EVAL_73 = _EVAL_455 & _EVAL_446;
  assign _EVAL_388 = _EVAL_220 & _EVAL_73;
  assign _EVAL_177 = _EVAL_145 & _EVAL_388;
  assign _EVAL_333 = _EVAL | _EVAL_314;
  assign _EVAL_328 = _EVAL_333 ? _EVAL_10 : _EVAL_23;
  assign _EVAL_204 = 8'h1 << _EVAL_328;
  assign _EVAL_82 = _EVAL_204[1];
  assign _EVAL_395 = _EVAL_333 ? _EVAL_9 : 1'h1;
  assign _EVAL_424 = _EVAL_82 & _EVAL_395;
  assign _EVAL_307 = _EVAL_333 ? _EVAL : _EVAL_48;
  assign _EVAL_240 = _EVAL_19 & _EVAL_307;
  assign _EVAL_429 = _EVAL_424 & _EVAL_240;
  assign _EVAL_410 = _EVAL_386[5];
  assign _EVAL_87 = _EVAL_410 & _EVAL_388;
  assign _EVAL_302 = _EVAL_286 - 4'h1;
  assign _EVAL_353 = _EVAL_204[3];
  assign _EVAL_110 = _EVAL_353 & _EVAL_395;
  assign _EVAL_329 = _EVAL_110 & _EVAL_240;
  assign _EVAL_129 = _EVAL_204[5];
  assign _EVAL_88 = _EVAL_129 & _EVAL_395;
  assign _EVAL_408 = _EVAL_333 == 1'h0;
  assign _EVAL_81 = _EVAL_19 & _EVAL;
  assign _EVAL_458 = _EVAL_386[3];
  assign _EVAL_253 = _EVAL_458 & _EVAL_388;
  assign _EVAL_357 = {{3'd0}, _EVAL_253};
  assign _EVAL_390 = _EVAL_386[4];
  assign _EVAL_243 = _EVAL_390 & _EVAL_388;
  assign _EVAL_407 = _EVAL_204[4];
  assign _EVAL_415 = _EVAL_407 & _EVAL_395;
  assign _EVAL_108 = _EVAL_415 & _EVAL_240;
  assign _EVAL_263 = _EVAL_364 | _EVAL_220;
  assign _EVAL_293 = _EVAL_263 & _EVAL_211;
  assign _EVAL_366 = 13'h3f << _EVAL_58;
  assign _EVAL_283 = _EVAL_315 ? _EVAL_293 : _EVAL_220;
  assign _EVAL_360 = _EVAL_141 & _EVAL_283;
  assign _EVAL_160 = _EVAL_204[2];
  assign _EVAL_294 = _EVAL_160 & _EVAL_395;
  assign _EVAL_139 = _EVAL_294 & _EVAL_240;
  assign _EVAL_351 = _EVAL_4 == 2'h3;
  assign _EVAL_191 = _EVAL_309 ? _EVAL_351 : _EVAL_426;
  assign _EVAL_439 = _EVAL_165 & _EVAL_388;
  assign _EVAL_275 = {{3'd0}, _EVAL_41};
  assign _EVAL_111 = _EVAL_386[2];
  assign _EVAL_152 = _EVAL_111 & _EVAL_388;
  assign _EVAL_133 = {{3'd0}, _EVAL_329};
  assign _EVAL_206 = _EVAL_286 == 4'h1;
  assign _EVAL_254 = _EVAL_366[5:0];
  assign _EVAL_393 = ~ _EVAL_254;
  assign _EVAL_62 = _EVAL_393[5:2];
  assign _EVAL_76 = _EVAL_315 ? _EVAL_62 : 4'h0;
  assign _EVAL_136 = _EVAL_76 == 4'h0;
  assign _EVAL_146 = _EVAL_206 | _EVAL_136;
  assign _EVAL_251 = _EVAL_146 == 1'h0;
  assign _EVAL_334 = _EVAL_386[7];
  assign _EVAL_181 = _EVAL_334 & _EVAL_388;
  assign _EVAL_227 = _EVAL_103 + _EVAL_181;
  assign _EVAL_277 = _EVAL_51[6:0];
  assign _EVAL_276 = _EVAL_128 + _EVAL_357;
  assign _EVAL_303 = _EVAL_276 - _EVAL_133;
  assign _EVAL_202 = _EVAL_204[6];
  assign _EVAL_134 = _EVAL_202 & _EVAL_395;
  assign _EVAL_77 = _EVAL_134 & _EVAL_240;
  assign _EVAL_392 = _EVAL_386[1];
  assign _EVAL_278 = _EVAL_392 & _EVAL_388;
  assign _EVAL_199 = {{3'd0}, _EVAL_108};
  assign _EVAL_385 = _EVAL_88 & _EVAL_240;
  assign _EVAL_449 = _EVAL_204[0];
  assign _EVAL_404 = _EVAL_449 & _EVAL_395;
  assign _EVAL_349 = _EVAL_404 & _EVAL_240;
  assign _EVAL_289 = _EVAL_204[7];
  assign _EVAL_313 = {{3'd0}, _EVAL_385};
  assign _EVAL_356 = {{3'd0}, _EVAL_87};
  assign _EVAL_384 = _EVAL_252 + _EVAL_356;
  assign _EVAL_300 = _EVAL_289 & _EVAL_395;
  assign _EVAL_322 = _EVAL_300 & _EVAL_240;
  assign _EVAL_311 = {{3'd0}, _EVAL_243};
  assign _EVAL_296 = _EVAL_158 + _EVAL_311;
  assign _EVAL_121 = 17'h3ff << _EVAL_58;
  assign _EVAL_282 = _EVAL_121[9:0];
  assign _EVAL_83 = ~ _EVAL_282;
  assign _EVAL_223 = {_EVAL_58, 7'h0};
  assign _EVAL_100 = _EVAL_275 | _EVAL_223;
  assign _EVAL_241 = Queue_1__EVAL_7;
  assign _EVAL_400 = _EVAL_9 == 1'h0;
  assign _EVAL_180 = {{3'd0}, _EVAL_177};
  assign _EVAL_427 = _EVAL_377 + _EVAL_180;
  assign _EVAL_236 = {{3'd0}, _EVAL_77};
  assign _EVAL_95 = {{2'd0}, _EVAL_152};
  assign _EVAL_431 = _EVAL_209 + _EVAL_95;
  assign _EVAL_394 = {{2'd0}, _EVAL_139};
  assign _EVAL_232 = _EVAL_431 - _EVAL_394;
  assign _EVAL_70 = _EVAL_241 == 1'h0;
  assign _EVAL_192 = _EVAL_212 + _EVAL_439;
  assign _EVAL_247 = _EVAL_4 != 2'h0;
  assign _EVAL_327 = _EVAL_247 | _EVAL_191;
  assign _EVAL_319 = _EVAL_360 & _EVAL_34;
  assign _EVAL_208 = _EVAL_22[9:7];
  assign _EVAL_147 = Queue_1__EVAL_13;
  assign _EVAL_92 = _EVAL_296 - _EVAL_199;
  assign _EVAL_285 = _EVAL_192 - _EVAL_349;
  assign _EVAL_389 = _EVAL_22[6:0];
  assign _EVAL_306 = _EVAL_58 >= 3'h2;
  assign _EVAL_423 = _EVAL_299 + _EVAL_278;
  assign _EVAL_85 = _EVAL_427 - _EVAL_236;
  assign _EVAL_79 = _EVAL_51[9:7];
  assign _EVAL_194 = _EVAL_227 - _EVAL_322;
  assign _EVAL_185 = _EVAL_455 & _EVAL_315;
  assign _EVAL_86 = _EVAL_16 != 2'h0;
  assign _EVAL_201 = _EVAL_384 - _EVAL_313;
  assign _EVAL_448 = _EVAL_423 - _EVAL_429;
  assign Queue__EVAL_0 = _EVAL_185 & _EVAL_263;
  assign Queue__EVAL_5 = _EVAL_54;
  assign _EVAL_26 = Queue__EVAL_10;
  assign _EVAL_24 = _EVAL_141 & _EVAL_283;
  assign Queue_1__EVAL_20 = _EVAL_241 ? _EVAL_27 : _EVAL_47;
  assign Queue_1__EVAL_18 = _EVAL_54;
  assign _EVAL_21 = Queue_1__EVAL_12;
  assign _EVAL_44 = Queue_1__EVAL_14;
  assign _EVAL_25 = _EVAL_333 ? _EVAL : _EVAL_48;
  assign Queue_1__EVAL_0 = _EVAL_43;
  assign _EVAL_37 = Queue_1__EVAL_8;
  assign _EVAL_55 = Queue_1__EVAL_12;
  assign _EVAL_0 = _EVAL_333 ? 3'h1 : 3'h0;
  assign _EVAL_18 = _EVAL_333 ? _EVAL_327 : 1'h0;
  assign Queue__EVAL_9 = _EVAL_15;
  assign Queue__EVAL_4 = _EVAL_59;
  assign _EVAL_28 = _EVAL_147 & _EVAL_70;
  assign Queue__EVAL_2 = _EVAL_206 | _EVAL_136;
  assign _EVAL_53 = _EVAL_19 & _EVAL_408;
  assign _EVAL_3 = Queue_1__EVAL_6;
  assign _EVAL_49 = Queue__EVAL_7;
  assign _EVAL_45 = Queue_1__EVAL_8;
  assign _EVAL_36 = _EVAL_333 ? _EVAL_208 : _EVAL_79;
  assign _EVAL_29 = Queue_1__EVAL;
  assign _EVAL_5 = Queue_1__EVAL_4;
  assign _EVAL_56 = Queue_1__EVAL;
  assign _EVAL_20 = Queue_1__EVAL_3;
  assign _EVAL_8 = _EVAL_333 ? _EVAL_191 : _EVAL_86;
  assign _EVAL_2 = _EVAL_19;
  assign _EVAL_50 = Queue_1__EVAL_10;
  assign Queue__EVAL_3 = _EVAL_32;
  assign Queue__EVAL_8 = _EVAL_11;
  assign Queue_1__EVAL_15 = _EVAL_306 ? 3'h2 : _EVAL_58;
  assign _EVAL_57 = Queue_1__EVAL_17;
  assign Queue_1__EVAL_21 = 7'h48 == _EVAL_41 ? 3'h0 : _EVAL_184;
  assign Queue_1__EVAL_11 = {{1'd0}, _EVAL_100};
  assign _EVAL_6 = Queue_1__EVAL_3;
  assign _EVAL_17 = Queue__EVAL_1;
  assign Queue_1__EVAL_5 = _EVAL_15;
  assign _EVAL_12 = _EVAL_333 ? _EVAL_389 : _EVAL_277;
  assign _EVAL_52 = Queue_1__EVAL_4;
  assign _EVAL_35 = _EVAL_38;
  assign _EVAL_42 = Queue_1__EVAL_14;
  assign _EVAL_46 = Queue_1__EVAL_16;
  assign _EVAL_14 = Queue_1__EVAL_16;
  assign Queue_1__EVAL_9 = _EVAL_434 == 1'h0;
  assign Queue_1__EVAL_19 = _EVAL_455 & _EVAL_446;
  assign _EVAL_1 = _EVAL_147 & _EVAL_241;
  assign Queue_1__EVAL_2 = _EVAL_83[9:2];
  assign _EVAL_30 = Queue_1__EVAL_6;
  assign _EVAL_31 = Queue__EVAL;
  assign _EVAL_40 = Queue_1__EVAL_10;
  assign _EVAL_33 = Queue_1__EVAL_17;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_89 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_103 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_128 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_148 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_158 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_196 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_209 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_212 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_252 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_286 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_299 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_309 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_314 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_364 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_377 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_398 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_426 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_430 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge _EVAL_54) begin
    if (_EVAL_152) begin
      _EVAL_89 <= _EVAL_315;
    end
    if (_EVAL_15) begin
      _EVAL_103 <= 1'h0;
    end else begin
      _EVAL_103 <= _EVAL_194;
    end
    if (_EVAL_15) begin
      _EVAL_128 <= 4'h0;
    end else begin
      _EVAL_128 <= _EVAL_303;
    end
    if (_EVAL_87) begin
      _EVAL_148 <= _EVAL_315;
    end
    if (_EVAL_15) begin
      _EVAL_158 <= 4'h0;
    end else begin
      _EVAL_158 <= _EVAL_92;
    end
    if (_EVAL_243) begin
      _EVAL_196 <= _EVAL_315;
    end
    if (_EVAL_15) begin
      _EVAL_209 <= 3'h0;
    end else begin
      _EVAL_209 <= _EVAL_232;
    end
    if (_EVAL_15) begin
      _EVAL_212 <= 1'h0;
    end else begin
      _EVAL_212 <= _EVAL_285;
    end
    if (_EVAL_15) begin
      _EVAL_252 <= 4'h0;
    end else begin
      _EVAL_252 <= _EVAL_201;
    end
    if (_EVAL_15) begin
      _EVAL_286 <= 4'h0;
    end else begin
      if (_EVAL_319) begin
        if (_EVAL_155) begin
          if (_EVAL_315) begin
            _EVAL_286 <= _EVAL_62;
          end else begin
            _EVAL_286 <= 4'h0;
          end
        end else begin
          _EVAL_286 <= _EVAL_302;
        end
      end
    end
    if (_EVAL_15) begin
      _EVAL_299 <= 1'h0;
    end else begin
      _EVAL_299 <= _EVAL_448;
    end
    if (_EVAL_15) begin
      _EVAL_309 <= 1'h1;
    end else begin
      if (_EVAL_81) begin
        _EVAL_309 <= _EVAL_9;
      end
    end
    if (_EVAL_15) begin
      _EVAL_314 <= 1'h0;
    end else begin
      if (_EVAL_81) begin
        _EVAL_314 <= _EVAL_400;
      end
    end
    if (_EVAL_15) begin
      _EVAL_364 <= 1'h0;
    end else begin
      if (_EVAL_319) begin
        _EVAL_364 <= _EVAL_251;
      end
    end
    if (_EVAL_15) begin
      _EVAL_377 <= 4'h0;
    end else begin
      _EVAL_377 <= _EVAL_85;
    end
    if (_EVAL_177) begin
      _EVAL_398 <= _EVAL_315;
    end
    if (_EVAL_309) begin
      _EVAL_426 <= _EVAL_351;
    end
    if (_EVAL_253) begin
      _EVAL_430 <= _EVAL_315;
    end
  end
endmodule
