//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
module SiFive__EVAL_74(
  output [5:0]  _EVAL,
  output        _EVAL_0,
  output [31:0] _EVAL_1,
  output [1:0]  _EVAL_2,
  output [2:0]  _EVAL_3,
  output [7:0]  _EVAL_4,
  output [31:0] _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  output        _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  output [1:0]  _EVAL_12,
  output [1:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [1:0]  _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [7:0]  _EVAL_17,
  input  [5:0]  _EVAL_18,
  output [31:0] _EVAL_19,
  input  [7:0]  _EVAL_20,
  output        _EVAL_21,
  input  [7:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [1:0]  _EVAL_28,
  input         _EVAL_29,
  output [7:0]  _EVAL_30,
  output [7:0]  _EVAL_31,
  input  [7:0]  _EVAL_32,
  input  [1:0]  _EVAL_33,
  input  [31:0] _EVAL_34,
  input  [31:0] _EVAL_35,
  input         _EVAL_36,
  input  [2:0]  _EVAL_37,
  input  [5:0]  _EVAL_38,
  output        _EVAL_39,
  output [7:0]  _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  output        _EVAL_44,
  output [1:0]  _EVAL_45,
  output [1:0]  _EVAL_46,
  input  [1:0]  _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  output [31:0] _EVAL_50,
  output        _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input  [31:0] _EVAL_54,
  output        _EVAL_55,
  output [5:0]  _EVAL_56,
  output        _EVAL_57,
  input         _EVAL_58,
  output [2:0]  _EVAL_59,
  output [1:0]  _EVAL_60
);
  assign _EVAL_13 = _EVAL_15;
  assign _EVAL_5 = _EVAL_35;
  assign _EVAL_1 = _EVAL_54;
  assign _EVAL_39 = _EVAL_24;
  assign _EVAL_9 = _EVAL_27;
  assign _EVAL_51 = _EVAL_42;
  assign _EVAL_40 = _EVAL_32;
  assign _EVAL_19 = _EVAL_14;
  assign _EVAL_25 = _EVAL_29;
  assign _EVAL_50 = _EVAL_34;
  assign _EVAL_30 = {_EVAL_38,_EVAL_33};
  assign _EVAL_43 = _EVAL_49;
  assign _EVAL_0 = _EVAL_53;
  assign _EVAL_3 = _EVAL_8;
  assign _EVAL = _EVAL_22[7:2];
  assign _EVAL_16 = _EVAL_11;
  assign _EVAL_41 = _EVAL_6;
  assign _EVAL_57 = _EVAL_36;
  assign _EVAL_56 = _EVAL_20[7:2];
  assign _EVAL_55 = _EVAL_26;
  assign _EVAL_21 = _EVAL_52;
  assign _EVAL_46 = _EVAL_22[1:0];
  assign _EVAL_48 = _EVAL_58;
  assign _EVAL_59 = _EVAL_37;
  assign _EVAL_45 = _EVAL_20[1:0];
  assign _EVAL_60 = _EVAL_47;
  assign _EVAL_2 = _EVAL_28;
  assign _EVAL_12 = _EVAL_7;
  assign _EVAL_44 = _EVAL_23;
  assign _EVAL_31 = {_EVAL_18,_EVAL_10};
  assign _EVAL_4 = _EVAL_17;
endmodule
