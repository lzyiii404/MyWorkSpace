//
// Copyright (c) 2016-2019 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000, 00000000-0000-0000-0000-0000000000000
//VCS coverage exclude_file
module SiFive_TLTestIndicator_assert(
  input         clock,
  input         reset,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [1:0]  auto_in_a_bits_size,
  input  [11:0] auto_in_a_bits_source,
  input  [14:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
  input         auto_in_d_ready,
  input  [13:0] _T_20_bits_extra,
  input         _T_20_bits_read,
  input         Queue__EVAL_1,
  input         Queue__EVAL_4
);
  wire  TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire [1:0] TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire [3:0] TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [14:0] TLMonitor__EVAL_7;
  wire [2:0] TLMonitor__EVAL_8;
  wire [2:0] TLMonitor__EVAL_9;
  wire [2:0] TLMonitor__EVAL_10;
  wire [1:0] TLMonitor__EVAL_11;
  wire [11:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [11:0] TLMonitor__EVAL_14;
  SiFive__EVAL_314_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  assign TLMonitor__EVAL_3 = clock;
  assign TLMonitor__EVAL_13 = reset;
  assign TLMonitor__EVAL_0 = Queue__EVAL_1;
  assign TLMonitor__EVAL = auto_in_a_valid;
  assign TLMonitor__EVAL_8 = auto_in_a_bits_opcode;
  assign TLMonitor__EVAL_10 = auto_in_a_bits_param;
  assign TLMonitor__EVAL_11 = auto_in_a_bits_size;
  assign TLMonitor__EVAL_12 = auto_in_a_bits_source;
  assign TLMonitor__EVAL_7 = auto_in_a_bits_address;
  assign TLMonitor__EVAL_5 = auto_in_a_bits_mask;
  assign TLMonitor__EVAL_4 = auto_in_a_bits_corrupt;
  assign TLMonitor__EVAL_6 = auto_in_d_ready;
  assign TLMonitor__EVAL_1 = Queue__EVAL_4;
  assign TLMonitor__EVAL_9 = {{2'd0}, _T_20_bits_read};
  assign TLMonitor__EVAL_2 = _T_20_bits_extra[1:0];
  assign TLMonitor__EVAL_14 = _T_20_bits_extra[13:2];

endmodule
